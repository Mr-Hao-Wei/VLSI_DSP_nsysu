`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// IIR Chebyshev bandstop filter testbench
// Structure: IIR Cascaded Second-Order Sections Direct Form II
// Total order: 6
// Cut-off freq.: 60 Hz
// Sampling freq.: 360 Hz
//
// Author: Abbiter Liu
//////////////////////////////////////////////////////////////////////////////////

module testbench_pli;

    reg clk;
    reg reset;
    reg signed [27:0] x;
    wire signed [27:0] y;

    // Instantiate the test filter
    chebyshev_bs_iir #(.WL(28)) u0 (
        .clk(clk), 
        .reset(reset),
        .x(x), 
        .y(y)
    );

    // Generate clock with 100ns period
    initial clk = 0;
    always #50 clk = ~clk;


    integer  ii;

    // Initialize and pass sinusoidal input data of 60Hz with sampling frequency of 360Hz   
    initial begin
        x = 0; reset = 1; clk = 0; 
        #100 reset = 1; 
        #200 reset = 0;
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111111110000000000000};
            #100 x={28'b0000010000110001000000000000};
            #100 x={28'b0000010001101010000000000000};
            #100 x={28'b0000010010101010000000000000};
            #100 x={28'b0000010011011001000000000000};
            #100 x={28'b0000010011010101000000000000};
            #100 x={28'b0000010010100011000000000000};
            #100 x={28'b0000010001100000000000000000};
            #100 x={28'b0000010000101010000000000000};
            #100 x={28'b0000001111111110000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000001111101011000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111101111000000000000};
            #100 x={28'b0000010000011011000000000000};
            #100 x={28'b0000010001001101000000000000};
            #100 x={28'b0000010010001010000000000000};
            #100 x={28'b0000010010111101000000000000};
            #100 x={28'b0000010011001100000000000000};
            #100 x={28'b0000010010110010000000000000};
            #100 x={28'b0000010001111001000000000000};
            #100 x={28'b0000010001000101000000000000};
            #100 x={28'b0000010000010111000000000000};
            #100 x={28'b0000001111110101000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111101011000000000000};
            #100 x={28'b0000001111101100000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000010000001101000000000000};
            #100 x={28'b0000010000111011000000000000};
            #100 x={28'b0000010001101100000000000000};
            #100 x={28'b0000010010101000000000000000};
            #100 x={28'b0000010011011001000000000000};
            #100 x={28'b0000010011101001000000000000};
            #100 x={28'b0000010011010000000000000000};
            #100 x={28'b0000010010011001000000000000};
            #100 x={28'b0000010001100000000000000000};
            #100 x={28'b0000010000101100000000000000};
            #100 x={28'b0000010000000011000000000000};
            #100 x={28'b0000001111110000000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111111011000000000000};
            #100 x={28'b0000010000101001000000000000};
            #100 x={28'b0000010001011100000000000000};
            #100 x={28'b0000010010001111000000000000};
            #100 x={28'b0000010011000011000000000000};
            #100 x={28'b0000010011011011000000000000};
            #100 x={28'b0000010011001010000000000000};
            #100 x={28'b0000010010010111000000000000};
            #100 x={28'b0000010001011100000000000000};
            #100 x={28'b0000010000100110000000000000};
            #100 x={28'b0000001111110110000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110011101000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110011101000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111110111000000000000};
            #100 x={28'b0000010000100100000000000000};
            #100 x={28'b0000010001010110000000000000};
            #100 x={28'b0000010010010000000000000000};
            #100 x={28'b0000010011000100000000000000};
            #100 x={28'b0000010011011100000000000000};
            #100 x={28'b0000010011010000000000000000};
            #100 x={28'b0000010010011110000000000000};
            #100 x={28'b0000010001100000000000000000};
            #100 x={28'b0000010000100011000000000000};
            #100 x={28'b0000001111110001000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110011010000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110011001000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110011101000000000000};
            #100 x={28'b0000001110011010000000000000};
            #100 x={28'b0000001110010111000000000000};
            #100 x={28'b0000001110011010000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110011101000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000010000001111000000000000};
            #100 x={28'b0000010000110111000000000000};
            #100 x={28'b0000010001100111000000000000};
            #100 x={28'b0000010010011101000000000000};
            #100 x={28'b0000010011000011000000000000};
            #100 x={28'b0000010011001000000000000000};
            #100 x={28'b0000010010100100000000000000};
            #100 x={28'b0000010001101010000000000000};
            #100 x={28'b0000010000110101000000000000};
            #100 x={28'b0000010000000000000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110011101000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110011001000000000000};
            #100 x={28'b0000001110011001000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110011010000000000000};
            #100 x={28'b0000001110011000000000000000};
            #100 x={28'b0000001110011000000000000000};
            #100 x={28'b0000001110011010000000000000};
            #100 x={28'b0000001110011101000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110011001000000000000};
            #100 x={28'b0000001110011001000000000000};
            #100 x={28'b0000001110011000000000000000};
            #100 x={28'b0000001110011000000000000000};
            #100 x={28'b0000001110011000000000000000};
            #100 x={28'b0000001110010111000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110011001000000000000};
            #100 x={28'b0000001110011001000000000000};
            #100 x={28'b0000001110010101000000000000};
            #100 x={28'b0000001110011010000000000000};
            #100 x={28'b0000001110011001000000000000};
            #100 x={28'b0000001110011001000000000000};
            #100 x={28'b0000001110010100000000000000};
            #100 x={28'b0000001110010011000000000000};
            #100 x={28'b0000001110011000000000000000};
            #100 x={28'b0000001110011010000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011101000000000000};
            #100 x={28'b0000001110011010000000000000};
            #100 x={28'b0000001110010111000000000000};
            #100 x={28'b0000001110011010000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110011101000000000000};
            #100 x={28'b0000001110011010000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011101000000000000};
            #100 x={28'b0000001110011101000000000000};
            #100 x={28'b0000001110011101000000000000};
            #100 x={28'b0000001110011101000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110011101000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110010010000000000000};
            #100 x={28'b0000001110010010000000000000};
            #100 x={28'b0000001110010101000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110011010000000000000};
            #100 x={28'b0000001110010101000000000000};
            #100 x={28'b0000001110010011000000000000};
            #100 x={28'b0000001110011000000000000000};
            #100 x={28'b0000001110010111000000000000};
            #100 x={28'b0000001110010111000000000000};
            #100 x={28'b0000001110010100000000000000};
            #100 x={28'b0000001110010101000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111110000000000000000};
            #100 x={28'b0000010000100101000000000000};
            #100 x={28'b0000010001011111000000000000};
            #100 x={28'b0000010010011100000000000000};
            #100 x={28'b0000010011001101000000000000};
            #100 x={28'b0000010011010101000000000000};
            #100 x={28'b0000010010101010000000000000};
            #100 x={28'b0000010001100111000000000000};
            #100 x={28'b0000010000101001000000000000};
            #100 x={28'b0000001111101101000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110010100000000000000};
            #100 x={28'b0000001110001111000000000000};
            #100 x={28'b0000001110001010000000000000};
            #100 x={28'b0000001110001101000000000000};
            #100 x={28'b0000001110010001000000000000};
            #100 x={28'b0000001110010001000000000000};
            #100 x={28'b0000001110010000000000000000};
            #100 x={28'b0000001110001111000000000000};
            #100 x={28'b0000001110001011000000000000};
            #100 x={28'b0000001110001101000000000000};
            #100 x={28'b0000001110001111000000000000};
            #100 x={28'b0000001110001110000000000000};
            #100 x={28'b0000001110010000000000000000};
            #100 x={28'b0000001110001111000000000000};
            #100 x={28'b0000001110001110000000000000};
            #100 x={28'b0000001110001110000000000000};
            #100 x={28'b0000001110010000000000000000};
            #100 x={28'b0000001110010010000000000000};
            #100 x={28'b0000001110001110000000000000};
            #100 x={28'b0000001110010000000000000000};
            #100 x={28'b0000001110001100000000000000};
            #100 x={28'b0000001110001110000000000000};
            #100 x={28'b0000001110001101000000000000};
            #100 x={28'b0000001110001111000000000000};
            #100 x={28'b0000001110001101000000000000};
            #100 x={28'b0000001110001110000000000000};
            #100 x={28'b0000001110001110000000000000};
            #100 x={28'b0000001110001100000000000000};
            #100 x={28'b0000001110001110000000000000};
            #100 x={28'b0000001110010000000000000000};
            #100 x={28'b0000001110001111000000000000};
            #100 x={28'b0000001110010000000000000000};
            #100 x={28'b0000001110001111000000000000};
            #100 x={28'b0000001110010001000000000000};
            #100 x={28'b0000001110010001000000000000};
            #100 x={28'b0000001110001111000000000000};
            #100 x={28'b0000001110010001000000000000};
            #100 x={28'b0000001110010000000000000000};
            #100 x={28'b0000001110001101000000000000};
            #100 x={28'b0000001110001111000000000000};
            #100 x={28'b0000001110010010000000000000};
            #100 x={28'b0000001110010100000000000000};
            #100 x={28'b0000001110010110000000000000};
            #100 x={28'b0000001110010100000000000000};
            #100 x={28'b0000001110001110000000000000};
            #100 x={28'b0000001110001110000000000000};
            #100 x={28'b0000001110001111000000000000};
            #100 x={28'b0000001110001111000000000000};
            #100 x={28'b0000001110010001000000000000};
            #100 x={28'b0000001110010001000000000000};
            #100 x={28'b0000001110010001000000000000};
            #100 x={28'b0000001110010110000000000000};
            #100 x={28'b0000001110011000000000000000};
            #100 x={28'b0000001110010111000000000000};
            #100 x={28'b0000001110010111000000000000};
            #100 x={28'b0000001110010101000000000000};
            #100 x={28'b0000001110010110000000000000};
            #100 x={28'b0000001110011000000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110011001000000000000};
            #100 x={28'b0000001110010111000000000000};
            #100 x={28'b0000001110010111000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000010000000010000000000000};
            #100 x={28'b0000010001000000000000000000};
            #100 x={28'b0000010010001011000000000000};
            #100 x={28'b0000010011011011000000000000};
            #100 x={28'b0000010100010001000000000000};
            #100 x={28'b0000010100010011000000000000};
            #100 x={28'b0000010011100010000000000000};
            #100 x={28'b0000010010010110000000000000};
            #100 x={28'b0000010001001110000000000000};
            #100 x={28'b0000010000011000000000000000};
            #100 x={28'b0000001111111101000000000000};
            #100 x={28'b0000001111110011000000000000};
            #100 x={28'b0000001111101100000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111101011000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000001111110000000000000000};
            #100 x={28'b0000001111110000000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000001111110011000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000001111101100000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000010000000011000000000000};
            #100 x={28'b0000010001000000000000000000};
            #100 x={28'b0000010010001011000000000000};
            #100 x={28'b0000010011010111000000000000};
            #100 x={28'b0000010100001001000000000000};
            #100 x={28'b0000010100000101000000000000};
            #100 x={28'b0000010011010001000000000000};
            #100 x={28'b0000010010001010000000000000};
            #100 x={28'b0000010001001000000000000000};
            #100 x={28'b0000010000010101000000000000};
            #100 x={28'b0000001111111100000000000000};
            #100 x={28'b0000001111110101000000000000};
            #100 x={28'b0000001111101101000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110011101000000000000};
            #100 x={28'b0000001110011101000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000010000010000000000000000};
            #100 x={28'b0000010001000110000000000000};
            #100 x={28'b0000010010000011000000000000};
            #100 x={28'b0000010011000011000000000000};
            #100 x={28'b0000010011110010000000000000};
            #100 x={28'b0000010011110100000000000000};
            #100 x={28'b0000010011000111000000000000};
            #100 x={28'b0000010010000110000000000000};
            #100 x={28'b0000010001000011000000000000};
            #100 x={28'b0000010000001001000000000000};
            #100 x={28'b0000001111101011000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111101011000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111101011000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000010000001110000000000000};
            #100 x={28'b0000010000111010000000000000};
            #100 x={28'b0000010001101101000000000000};
            #100 x={28'b0000010010100110000000000000};
            #100 x={28'b0000010011010100000000000000};
            #100 x={28'b0000010011100101000000000000};
            #100 x={28'b0000010011001011000000000000};
            #100 x={28'b0000010010010011000000000000};
            #100 x={28'b0000010001010101000000000000};
            #100 x={28'b0000010000100001000000000000};
            #100 x={28'b0000001111111000000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111110000000000000000};
            #100 x={28'b0000010000011111000000000000};
            #100 x={28'b0000010001010101000000000000};
            #100 x={28'b0000010010010101000000000000};
            #100 x={28'b0000010011001110000000000000};
            #100 x={28'b0000010011101001000000000000};
            #100 x={28'b0000010011011001000000000000};
            #100 x={28'b0000010010101010000000000000};
            #100 x={28'b0000010001110010000000000000};
            #100 x={28'b0000010000111100000000000000};
            #100 x={28'b0000010000000110000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111111000000000000000};
            #100 x={28'b0000010000100110000000000000};
            #100 x={28'b0000010001100000000000000000};
            #100 x={28'b0000010010100010000000000000};
            #100 x={28'b0000010011011011000000000000};
            #100 x={28'b0000010011101110000000000000};
            #100 x={28'b0000010011001111000000000000};
            #100 x={28'b0000010010010011000000000000};
            #100 x={28'b0000010001011010000000000000};
            #100 x={28'b0000010000100100000000000000};
            #100 x={28'b0000001111111101000000000000};
            #100 x={28'b0000001111101101000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111101011000000000000};
            #100 x={28'b0000001111101011000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111101100000000000000};
            #100 x={28'b0000001111101011000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000001111101011000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000010000000110000000000000};
            #100 x={28'b0000010000111001000000000000};
            #100 x={28'b0000010001111000000000000000};
            #100 x={28'b0000010010111110000000000000};
            #100 x={28'b0000010011101110000000000000};
            #100 x={28'b0000010011110011000000000000};
            #100 x={28'b0000010011000111000000000000};
            #100 x={28'b0000010010000110000000000000};
            #100 x={28'b0000010001001011000000000000};
            #100 x={28'b0000010000100010000000000000};
            #100 x={28'b0000010000001011000000000000};
            #100 x={28'b0000010000000100000000000000};
            #100 x={28'b0000010000000001000000000000};
            #100 x={28'b0000001111111011000000000000};
            #100 x={28'b0000001111110110000000000000};
            #100 x={28'b0000001111110010000000000000};
            #100 x={28'b0000001111101011000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111101100000000000000};
            #100 x={28'b0000001111101111000000000000};
            #100 x={28'b0000001111101111000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000001111110001000000000000};
            #100 x={28'b0000001111110100000000000000};
            #100 x={28'b0000001111110110000000000000};
            #100 x={28'b0000001111110011000000000000};
            #100 x={28'b0000001111101111000000000000};
            #100 x={28'b0000001111110010000000000000};
            #100 x={28'b0000001111110101000000000000};
            #100 x={28'b0000001111110010000000000000};
            #100 x={28'b0000001111110001000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000001111101011000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111101100000000000000};
            #100 x={28'b0000001111110100000000000000};
            #100 x={28'b0000001111111000000000000000};
            #100 x={28'b0000001111110100000000000000};
            #100 x={28'b0000001111110000000000000000};
            #100 x={28'b0000001111101101000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000001111101111000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111110111000000000000};
            #100 x={28'b0000010000100101000000000000};
            #100 x={28'b0000010001011101000000000000};
            #100 x={28'b0000010010011111000000000000};
            #100 x={28'b0000010011011001000000000000};
            #100 x={28'b0000010011100111000000000000};
            #100 x={28'b0000010011000111000000000000};
            #100 x={28'b0000010010001101000000000000};
            #100 x={28'b0000010001001111000000000000};
            #100 x={28'b0000010000011110000000000000};
            #100 x={28'b0000010000001010000000000000};
            #100 x={28'b0000010000001011000000000000};
            #100 x={28'b0000010000000111000000000000};
            #100 x={28'b0000010000000000000000000000};
            #100 x={28'b0000001111110100000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111101100000000000000};
            #100 x={28'b0000001111101100000000000000};
            #100 x={28'b0000001111101011000000000000};
            #100 x={28'b0000001111101011000000000000};
            #100 x={28'b0000001111101011000000000000};
            #100 x={28'b0000001111101100000000000000};
            #100 x={28'b0000001111101111000000000000};
            #100 x={28'b0000001111110000000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000001111101100000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111101011000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111101100000000000000};
            #100 x={28'b0000001111101011000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111110001000000000000};
            #100 x={28'b0000010000010101000000000000};
            #100 x={28'b0000010001000011000000000000};
            #100 x={28'b0000010001111111000000000000};
            #100 x={28'b0000010010110011000000000000};
            #100 x={28'b0000010010111110000000000000};
            #100 x={28'b0000010010010111000000000000};
            #100 x={28'b0000010001010110000000000000};
            #100 x={28'b0000010000011110000000000000};
            #100 x={28'b0000001111110111000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110011101000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110011010000000000000};
            #100 x={28'b0000001110010110000000000000};
            #100 x={28'b0000001110011000000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110011010000000000000};
            #100 x={28'b0000001110011000000000000000};
            #100 x={28'b0000001110011001000000000000};
            #100 x={28'b0000001110011000000000000000};
            #100 x={28'b0000001110010101000000000000};
            #100 x={28'b0000001110010111000000000000};
            #100 x={28'b0000001110011000000000000000};
            #100 x={28'b0000001110011000000000000000};
            #100 x={28'b0000001110010111000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011010000000000000};
            #100 x={28'b0000001110010010000000000000};
            #100 x={28'b0000001110001111000000000000};
            #100 x={28'b0000001110010010000000000000};
            #100 x={28'b0000001110010111000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110011001000000000000};
            #100 x={28'b0000001110010111000000000000};
            #100 x={28'b0000001110010111000000000000};
            #100 x={28'b0000001110011000000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110011101000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000001111101101000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111111101000000000000};
            #100 x={28'b0000010000101100000000000000};
            #100 x={28'b0000010001100010000000000000};
            #100 x={28'b0000010010100010000000000000};
            #100 x={28'b0000010011011100000000000000};
            #100 x={28'b0000010011111010000000000000};
            #100 x={28'b0000010011100111000000000000};
            #100 x={28'b0000010010110010000000000000};
            #100 x={28'b0000010001111001000000000000};
            #100 x={28'b0000010001000101000000000000};
            #100 x={28'b0000010000011010000000000000};
            #100 x={28'b0000010000001001000000000000};
            #100 x={28'b0000010000001000000000000000};
            #100 x={28'b0000010000000010000000000000};
            #100 x={28'b0000001111111000000000000000};
            #100 x={28'b0000001111101111000000000000};
            #100 x={28'b0000001111101101000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111101101000000000000};
            #100 x={28'b0000001111101111000000000000};
            #100 x={28'b0000001111110000000000000000};
            #100 x={28'b0000001111110010000000000000};
            #100 x={28'b0000001111110011000000000000};
            #100 x={28'b0000001111110010000000000000};
            #100 x={28'b0000001111110010000000000000};
            #100 x={28'b0000001111110010000000000000};
            #100 x={28'b0000001111110011000000000000};
            #100 x={28'b0000001111110010000000000000};
            #100 x={28'b0000001111110100000000000000};
            #100 x={28'b0000001111110110000000000000};
            #100 x={28'b0000001111111000000000000000};
            #100 x={28'b0000001111111000000000000000};
            #100 x={28'b0000001111110010000000000000};
            #100 x={28'b0000001111110001000000000000};
            #100 x={28'b0000001111110000000000000000};
            #100 x={28'b0000001111110010000000000000};
            #100 x={28'b0000001111110001000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000001111101111000000000000};
            #100 x={28'b0000001111101100000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111111101000000000000};
            #100 x={28'b0000010000101110000000000000};
            #100 x={28'b0000010001100011000000000000};
            #100 x={28'b0000010010100010000000000000};
            #100 x={28'b0000010011010110000000000000};
            #100 x={28'b0000010011101100000000000000};
            #100 x={28'b0000010011010000000000000000};
            #100 x={28'b0000010010011011000000000000};
            #100 x={28'b0000010001100101000000000000};
            #100 x={28'b0000010000110101000000000000};
            #100 x={28'b0000010000001111000000000000};
            #100 x={28'b0000010000000010000000000000};
            #100 x={28'b0000010000000000000000000000};
            #100 x={28'b0000001111111011000000000000};
            #100 x={28'b0000001111110100000000000000};
            #100 x={28'b0000001111101100000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111101011000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000010000001111000000000000};
            #100 x={28'b0000010000111111000000000000};
            #100 x={28'b0000010001111100000000000000};
            #100 x={28'b0000010010101101000000000000};
            #100 x={28'b0000010010111100000000000000};
            #100 x={28'b0000010010011101000000000000};
            #100 x={28'b0000010001101100000000000000};
            #100 x={28'b0000010000111100000000000000};
            #100 x={28'b0000010000010010000000000000};
            #100 x={28'b0000001111101100000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110010110000000000000};
            #100 x={28'b0000001110010101000000000000};
            #100 x={28'b0000001110011001000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110011001000000000000};
            #100 x={28'b0000001110010101000000000000};
            #100 x={28'b0000001110010000000000000000};
            #100 x={28'b0000001110010010000000000000};
            #100 x={28'b0000001110010101000000000000};
            #100 x={28'b0000001110011001000000000000};
            #100 x={28'b0000001110010110000000000000};
            #100 x={28'b0000001110010011000000000000};
            #100 x={28'b0000001110010001000000000000};
            #100 x={28'b0000001110010001000000000000};
            #100 x={28'b0000001110010100000000000000};
            #100 x={28'b0000001110010011000000000000};
            #100 x={28'b0000001110010101000000000000};
            #100 x={28'b0000001110010101000000000000};
            #100 x={28'b0000001110010100000000000000};
            #100 x={28'b0000001110010001000000000000};
            #100 x={28'b0000001110010100000000000000};
            #100 x={28'b0000001110010100000000000000};
            #100 x={28'b0000001110011000000000000000};
            #100 x={28'b0000001110010111000000000000};
            #100 x={28'b0000001110010010000000000000};
            #100 x={28'b0000001110010001000000000000};
            #100 x={28'b0000001110010010000000000000};
            #100 x={28'b0000001110010110000000000000};
            #100 x={28'b0000001110011000000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110011000000000000000};
            #100 x={28'b0000001110010010000000000000};
            #100 x={28'b0000001110010000000000000000};
            #100 x={28'b0000001110010011000000000000};
            #100 x={28'b0000001110010110000000000000};
            #100 x={28'b0000001110010101000000000000};
            #100 x={28'b0000001110010101000000000000};
            #100 x={28'b0000001110010010000000000000};
            #100 x={28'b0000001110010001000000000000};
            #100 x={28'b0000001110010100000000000000};
            #100 x={28'b0000001110010100000000000000};
            #100 x={28'b0000001110010100000000000000};
            #100 x={28'b0000001110010011000000000000};
            #100 x={28'b0000001110010010000000000000};
            #100 x={28'b0000001110010101000000000000};
            #100 x={28'b0000001110010110000000000000};
            #100 x={28'b0000001110010111000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110010111000000000000};
            #100 x={28'b0000001110010001000000000000};
            #100 x={28'b0000001110010100000000000000};
            #100 x={28'b0000001110011010000000000000};
            #100 x={28'b0000001110011101000000000000};
            #100 x={28'b0000001110010111000000000000};
            #100 x={28'b0000001110011000000000000000};
            #100 x={28'b0000001110011001000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110011101000000000000};
            #100 x={28'b0000001110011101000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000010000010100000000000000};
            #100 x={28'b0000010001000011000000000000};
            #100 x={28'b0000010001111110000000000000};
            #100 x={28'b0000010010111100000000000000};
            #100 x={28'b0000010011100011000000000000};
            #100 x={28'b0000010011011110000000000000};
            #100 x={28'b0000010010110100000000000000};
            #100 x={28'b0000010001111110000000000000};
            #100 x={28'b0000010001001101000000000000};
            #100 x={28'b0000010000100000000000000000};
            #100 x={28'b0000010000000100000000000000};
            #100 x={28'b0000001111111101000000000000};
            #100 x={28'b0000001111111010000000000000};
            #100 x={28'b0000001111110001000000000000};
            #100 x={28'b0000001111101011000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000001111110001000000000000};
            #100 x={28'b0000001111110100000000000000};
            #100 x={28'b0000001111110110000000000000};
            #100 x={28'b0000001111110010000000000000};
            #100 x={28'b0000001111110011000000000000};
            #100 x={28'b0000001111110101000000000000};
            #100 x={28'b0000001111110111000000000000};
            #100 x={28'b0000001111111010000000000000};
            #100 x={28'b0000001111111010000000000000};
            #100 x={28'b0000001111111001000000000000};
            #100 x={28'b0000001111111000000000000000};
            #100 x={28'b0000001111111010000000000000};
            #100 x={28'b0000001111111010000000000000};
            #100 x={28'b0000001111111010000000000000};
            #100 x={28'b0000001111111001000000000000};
            #100 x={28'b0000001111110011000000000000};
            #100 x={28'b0000001111110011000000000000};
            #100 x={28'b0000001111110100000000000000};
            #100 x={28'b0000001111110111000000000000};
            #100 x={28'b0000001111110110000000000000};
            #100 x={28'b0000001111110001000000000000};
            #100 x={28'b0000001111101100000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111110100000000000000};
            #100 x={28'b0000001111111010000000000000};
            #100 x={28'b0000001111111010000000000000};
            #100 x={28'b0000001111110100000000000000};
            #100 x={28'b0000001111101111000000000000};
            #100 x={28'b0000001111110000000000000000};
            #100 x={28'b0000001111110011000000000000};
            #100 x={28'b0000001111110001000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000001111101011000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000010000001010000000000000};
            #100 x={28'b0000010000111111000000000000};
            #100 x={28'b0000010001111110000000000000};
            #100 x={28'b0000010011000100000000000000};
            #100 x={28'b0000010011110010000000000000};
            #100 x={28'b0000010011110000000000000000};
            #100 x={28'b0000010010111000000000000000};
            #100 x={28'b0000010001111001000000000000};
            #100 x={28'b0000010001000111000000000000};
            #100 x={28'b0000010000011111000000000000};
            #100 x={28'b0000010000001111000000000000};
            #100 x={28'b0000010000001110000000000000};
            #100 x={28'b0000010000001010000000000000};
            #100 x={28'b0000010000000011000000000000};
            #100 x={28'b0000001111111101000000000000};
            #100 x={28'b0000001111110011000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111110000000000000000};
            #100 x={28'b0000001111110000000000000000};
            #100 x={28'b0000001111101111000000000000};
            #100 x={28'b0000001111101101000000000000};
            #100 x={28'b0000001111101101000000000000};
            #100 x={28'b0000001111110011000000000000};
            #100 x={28'b0000001111110100000000000000};
            #100 x={28'b0000001111110110000000000000};
            #100 x={28'b0000001111110111000000000000};
            #100 x={28'b0000001111110110000000000000};
            #100 x={28'b0000001111111001000000000000};
            #100 x={28'b0000001111111010000000000000};
            #100 x={28'b0000001111111000000000000000};
            #100 x={28'b0000001111111000000000000000};
            #100 x={28'b0000001111110110000000000000};
            #100 x={28'b0000001111110011000000000000};
            #100 x={28'b0000001111110001000000000000};
            #100 x={28'b0000001111110010000000000000};
            #100 x={28'b0000001111110100000000000000};
            #100 x={28'b0000001111110010000000000000};
            #100 x={28'b0000001111101111000000000000};
            #100 x={28'b0000001111101011000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111101011000000000000};
            #100 x={28'b0000001111110001000000000000};
            #100 x={28'b0000001111110011000000000000};
            #100 x={28'b0000001111101111000000000000};
            #100 x={28'b0000001111101011000000000000};
            #100 x={28'b0000001111101100000000000000};
            #100 x={28'b0000001111101101000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000010000001001000000000000};
            #100 x={28'b0000010000111000000000000000};
            #100 x={28'b0000010001110100000000000000};
            #100 x={28'b0000010010111000000000000000};
            #100 x={28'b0000010011101000000000000000};
            #100 x={28'b0000010011101100000000000000};
            #100 x={28'b0000010010111111000000000000};
            #100 x={28'b0000010010000010000000000000};
            #100 x={28'b0000010001001000000000000000};
            #100 x={28'b0000010000011011000000000000};
            #100 x={28'b0000010000000101000000000000};
            #100 x={28'b0000010000000101000000000000};
            #100 x={28'b0000010000000001000000000000};
            #100 x={28'b0000001111111101000000000000};
            #100 x={28'b0000001111110101000000000000};
            #100 x={28'b0000001111101100000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111101011000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111101011000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111101011000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000010000010001000000000000};
            #100 x={28'b0000010001000101000000000000};
            #100 x={28'b0000010010000011000000000000};
            #100 x={28'b0000010010111011000000000000};
            #100 x={28'b0000010011010100000000000000};
            #100 x={28'b0000010010111111000000000000};
            #100 x={28'b0000010010001000000000000000};
            #100 x={28'b0000010001001100000000000000};
            #100 x={28'b0000010000011000000000000000};
            #100 x={28'b0000001111110111000000000000};
            #100 x={28'b0000001111110000000000000000};
            #100 x={28'b0000001111101111000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111111111000000000000};
            #100 x={28'b0000010000101111000000000000};
            #100 x={28'b0000010001101110000000000000};
            #100 x={28'b0000010010101000000000000000};
            #100 x={28'b0000010010111110000000000000};
            #100 x={28'b0000010010101000000000000000};
            #100 x={28'b0000010001110001000000000000};
            #100 x={28'b0000010000111100000000000000};
            #100 x={28'b0000010000001111000000000000};
            #100 x={28'b0000001111101111000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110011000000000000000};
            #100 x={28'b0000001110011000000000000000};
            #100 x={28'b0000001110011000000000000000};
            #100 x={28'b0000001110011010000000000000};
            #100 x={28'b0000001110011010000000000000};
            #100 x={28'b0000001110011000000000000000};
            #100 x={28'b0000001110010111000000000000};
            #100 x={28'b0000001110010101000000000000};
            #100 x={28'b0000001110010111000000000000};
            #100 x={28'b0000001110011000000000000000};
            #100 x={28'b0000001110010111000000000000};
            #100 x={28'b0000001110010110000000000000};
            #100 x={28'b0000001110010101000000000000};
            #100 x={28'b0000001110010111000000000000};
            #100 x={28'b0000001110011001000000000000};
            #100 x={28'b0000001110011010000000000000};
            #100 x={28'b0000001110010111000000000000};
            #100 x={28'b0000001110010111000000000000};
            #100 x={28'b0000001110010110000000000000};
            #100 x={28'b0000001110011010000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110011001000000000000};
            #100 x={28'b0000001110011001000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011101000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111111110000000000000};
            #100 x={28'b0000010000101010000000000000};
            #100 x={28'b0000010001100011000000000000};
            #100 x={28'b0000010010100001000000000000};
            #100 x={28'b0000010011000110000000000000};
            #100 x={28'b0000010010110100000000000000};
            #100 x={28'b0000010001111011000000000000};
            #100 x={28'b0000010001000010000000000000};
            #100 x={28'b0000010000010011000000000000};
            #100 x={28'b0000001111111000000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110011101000000000000};
            #100 x={28'b0000001110011101000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011101000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110011101000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011101000000000000};
            #100 x={28'b0000001110011010000000000000};
            #100 x={28'b0000001110011101000000000000};
            #100 x={28'b0000001110011101000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110011101000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011101000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110011101000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110011101000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111110000000000000000};
            #100 x={28'b0000010000100000000000000000};
            #100 x={28'b0000010001100000000000000000};
            #100 x={28'b0000010010011100000000000000};
            #100 x={28'b0000010010110100000000000000};
            #100 x={28'b0000010010011011000000000000};
            #100 x={28'b0000010001011100000000000000};
            #100 x={28'b0000010000100110000000000000};
            #100 x={28'b0000001111110111000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110011010000000000000};
            #100 x={28'b0000001110011001000000000000};
            #100 x={28'b0000001110011000000000000000};
            #100 x={28'b0000001110011000000000000000};
            #100 x={28'b0000001110010110000000000000};
            #100 x={28'b0000001110010011000000000000};
            #100 x={28'b0000001110010011000000000000};
            #100 x={28'b0000001110010100000000000000};
            #100 x={28'b0000001110010101000000000000};
            #100 x={28'b0000001110010111000000000000};
            #100 x={28'b0000001110011001000000000000};
            #100 x={28'b0000001110011000000000000000};
            #100 x={28'b0000001110010101000000000000};
            #100 x={28'b0000001110010011000000000000};
            #100 x={28'b0000001110010101000000000000};
            #100 x={28'b0000001110011000000000000000};
            #100 x={28'b0000001110010110000000000000};
            #100 x={28'b0000001110010101000000000000};
            #100 x={28'b0000001110010100000000000000};
            #100 x={28'b0000001110010101000000000000};
            #100 x={28'b0000001110011000000000000000};
            #100 x={28'b0000001110011001000000000000};
            #100 x={28'b0000001110010100000000000000};
            #100 x={28'b0000001110010110000000000000};
            #100 x={28'b0000001110010011000000000000};
            #100 x={28'b0000001110010011000000000000};
            #100 x={28'b0000001110010110000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110011000000000000000};
            #100 x={28'b0000001110010010000000000000};
            #100 x={28'b0000001110010001000000000000};
            #100 x={28'b0000001110010110000000000000};
            #100 x={28'b0000001110011010000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110011000000000000000};
            #100 x={28'b0000001110010111000000000000};
            #100 x={28'b0000001110011000000000000000};
            #100 x={28'b0000001110011010000000000000};
            #100 x={28'b0000001110011010000000000000};
            #100 x={28'b0000001110011001000000000000};
            #100 x={28'b0000001110011010000000000000};
            #100 x={28'b0000001110011000000000000000};
            #100 x={28'b0000001110011000000000000000};
            #100 x={28'b0000001110011001000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011101000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011101000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011101000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111110000000000000000};
            #100 x={28'b0000010000101001000000000000};
            #100 x={28'b0000010001100110000000000000};
            #100 x={28'b0000010010101011000000000000};
            #100 x={28'b0000010011011100000000000000};
            #100 x={28'b0000010011011101000000000000};
            #100 x={28'b0000010010101111000000000000};
            #100 x={28'b0000010001110011000000000000};
            #100 x={28'b0000010000110010000000000000};
            #100 x={28'b0000001111111010000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110011000000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110011010000000000000};
            #100 x={28'b0000001110011001000000000000};
            #100 x={28'b0000001110010110000000000000};
            #100 x={28'b0000001110010110000000000000};
            #100 x={28'b0000001110011000000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110011010000000000000};
            #100 x={28'b0000001110011010000000000000};
            #100 x={28'b0000001110010101000000000000};
            #100 x={28'b0000001110010111000000000000};
            #100 x={28'b0000001110010111000000000000};
            #100 x={28'b0000001110011010000000000000};
            #100 x={28'b0000001110011001000000000000};
            #100 x={28'b0000001110010110000000000000};
            #100 x={28'b0000001110010110000000000000};
            #100 x={28'b0000001110010110000000000000};
            #100 x={28'b0000001110011001000000000000};
            #100 x={28'b0000001110011010000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110011010000000000000};
            #100 x={28'b0000001110011001000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110011101000000000000};
            #100 x={28'b0000001110011101000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111111010000000000000};
            #100 x={28'b0000010000101100000000000000};
            #100 x={28'b0000010001101001000000000000};
            #100 x={28'b0000010010101010000000000000};
            #100 x={28'b0000010011100101000000000000};
            #100 x={28'b0000010011111101000000000000};
            #100 x={28'b0000010011011100000000000000};
            #100 x={28'b0000010010100001000000000000};
            #100 x={28'b0000010001100011000000000000};
            #100 x={28'b0000010000101111000000000000};
            #100 x={28'b0000010000010001000000000000};
            #100 x={28'b0000010000001011000000000000};
            #100 x={28'b0000010000001001000000000000};
            #100 x={28'b0000001111111111000000000000};
            #100 x={28'b0000001111110110000000000000};
            #100 x={28'b0000001111101100000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111101100000000000000};
            #100 x={28'b0000001111101111000000000000};
            #100 x={28'b0000001111101111000000000000};
            #100 x={28'b0000001111101100000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111101101000000000000};
            #100 x={28'b0000001111101111000000000000};
            #100 x={28'b0000001111101100000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111101100000000000000};
            #100 x={28'b0000001111101011000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111101100000000000000};
            #100 x={28'b0000010000010111000000000000};
            #100 x={28'b0000010001000101000000000000};
            #100 x={28'b0000010001111110000000000000};
            #100 x={28'b0000010010111010000000000000};
            #100 x={28'b0000010011010111000000000000};
            #100 x={28'b0000010011000111000000000000};
            #100 x={28'b0000010010010010000000000000};
            #100 x={28'b0000010001011011000000000000};
            #100 x={28'b0000010000100101000000000000};
            #100 x={28'b0000010000000010000000000000};
            #100 x={28'b0000001111110110000000000000};
            #100 x={28'b0000001111110100000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110011101000000000000};
            #100 x={28'b0000001110011010000000000000};
            #100 x={28'b0000001110011101000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111101111000000000000};
            #100 x={28'b0000010000100001000000000000};
            #100 x={28'b0000010001011000000000000000};
            #100 x={28'b0000010010011101000000000000};
            #100 x={28'b0000010011010110000000000000};
            #100 x={28'b0000010011110000000000000000};
            #100 x={28'b0000010011011000000000000000};
            #100 x={28'b0000010010100000000000000000};
            #100 x={28'b0000010001100100000000000000};
            #100 x={28'b0000010000101111000000000000};
            #100 x={28'b0000010000001111000000000000};
            #100 x={28'b0000010000000011000000000000};
            #100 x={28'b0000010000000000000000000000};
            #100 x={28'b0000001111110111000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111101100000000000000};
            #100 x={28'b0000001111101111000000000000};
            #100 x={28'b0000001111110001000000000000};
            #100 x={28'b0000001111110001000000000000};
            #100 x={28'b0000001111101111000000000000};
            #100 x={28'b0000001111101111000000000000};
            #100 x={28'b0000001111110100000000000000};
            #100 x={28'b0000001111110110000000000000};
            #100 x={28'b0000001111111000000000000000};
            #100 x={28'b0000001111111010000000000000};
            #100 x={28'b0000001111111000000000000000};
            #100 x={28'b0000001111110110000000000000};
            #100 x={28'b0000001111111010000000000000};
            #100 x={28'b0000001111111011000000000000};
            #100 x={28'b0000001111111001000000000000};
            #100 x={28'b0000001111111001000000000000};
            #100 x={28'b0000001111110110000000000000};
            #100 x={28'b0000001111110101000000000000};
            #100 x={28'b0000001111110110000000000000};
            #100 x={28'b0000001111110011000000000000};
            #100 x={28'b0000001111110000000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000001111110010000000000000};
            #100 x={28'b0000001111110111000000000000};
            #100 x={28'b0000001111110101000000000000};
            #100 x={28'b0000001111110011000000000000};
            #100 x={28'b0000001111110001000000000000};
            #100 x={28'b0000001111101111000000000000};
            #100 x={28'b0000001111110011000000000000};
            #100 x={28'b0000001111110100000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111101100000000000000};
            #100 x={28'b0000001111101100000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000010000001011000000000000};
            #100 x={28'b0000010000111100000000000000};
            #100 x={28'b0000010001110010000000000000};
            #100 x={28'b0000010010101101000000000000};
            #100 x={28'b0000010011100011000000000000};
            #100 x={28'b0000010011110111000000000000};
            #100 x={28'b0000010011011000000000000000};
            #100 x={28'b0000010010011111000000000000};
            #100 x={28'b0000010001100111000000000000};
            #100 x={28'b0000010000110011000000000000};
            #100 x={28'b0000010000001101000000000000};
            #100 x={28'b0000010000000000000000000000};
            #100 x={28'b0000010000000000000000000000};
            #100 x={28'b0000001111111011000000000000};
            #100 x={28'b0000001111110100000000000000};
            #100 x={28'b0000001111101101000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111101100000000000000};
            #100 x={28'b0000001111110001000000000000};
            #100 x={28'b0000001111110001000000000000};
            #100 x={28'b0000001111110011000000000000};
            #100 x={28'b0000001111110010000000000000};
            #100 x={28'b0000001111110100000000000000};
            #100 x={28'b0000001111110111000000000000};
            #100 x={28'b0000001111111011000000000000};
            #100 x={28'b0000001111111011000000000000};
            #100 x={28'b0000001111111010000000000000};
            #100 x={28'b0000001111111001000000000000};
            #100 x={28'b0000001111111110000000000000};
            #100 x={28'b0000001111111110000000000000};
            #100 x={28'b0000010000000001000000000000};
            #100 x={28'b0000001111111111000000000000};
            #100 x={28'b0000010000000011000000000000};
            #100 x={28'b0000010000000101000000000000};
            #100 x={28'b0000010000001001000000000000};
            #100 x={28'b0000010000001011000000000000};
            #100 x={28'b0000010000001011000000000000};
            #100 x={28'b0000010000000111000000000000};
            #100 x={28'b0000010000000011000000000000};
            #100 x={28'b0000001111111111000000000000};
            #100 x={28'b0000010000000001000000000000};
            #100 x={28'b0000010000000010000000000000};
            #100 x={28'b0000010000000100000000000000};
            #100 x={28'b0000010000000101000000000000};
            #100 x={28'b0000010000000011000000000000};
            #100 x={28'b0000010000000010000000000000};
            #100 x={28'b0000001111111110000000000000};
            #100 x={28'b0000001111111000000000000000};
            #100 x={28'b0000001111110100000000000000};
            #100 x={28'b0000001111110000000000000000};
            #100 x={28'b0000001111101100000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000001111101111000000000000};
            #100 x={28'b0000001111101111000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000001111110001000000000000};
            #100 x={28'b0000001111110101000000000000};
            #100 x={28'b0000001111111010000000000000};
            #100 x={28'b0000001111111101000000000000};
            #100 x={28'b0000010000000011000000000000};
            #100 x={28'b0000010000000011000000000000};
            #100 x={28'b0000010000000001000000000000};
            #100 x={28'b0000001111111110000000000000};
            #100 x={28'b0000001111111110000000000000};
            #100 x={28'b0000001111111001000000000000};
            #100 x={28'b0000001111111000000000000000};
            #100 x={28'b0000001111110101000000000000};
            #100 x={28'b0000001111110110000000000000};
            #100 x={28'b0000001111110101000000000000};
            #100 x={28'b0000001111110100000000000000};
            #100 x={28'b0000001111110100000000000000};
            #100 x={28'b0000001111111000000000000000};
            #100 x={28'b0000001111111101000000000000};
            #100 x={28'b0000001111111001000000000000};
            #100 x={28'b0000001111110010000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000010000000000000000000000};
            #100 x={28'b0000010000101001000000000000};
            #100 x={28'b0000010001010111000000000000};
            #100 x={28'b0000010010001101000000000000};
            #100 x={28'b0000010011001010000000000000};
            #100 x={28'b0000010011110010000000000000};
            #100 x={28'b0000010011110100000000000000};
            #100 x={28'b0000010011001100000000000000};
            #100 x={28'b0000010010010110000000000000};
            #100 x={28'b0000010001100111000000000000};
            #100 x={28'b0000010000111001000000000000};
            #100 x={28'b0000010000010101000000000000};
            #100 x={28'b0000001111111111000000000000};
            #100 x={28'b0000001111111010000000000000};
            #100 x={28'b0000001111110100000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111110000000000000000};
            #100 x={28'b0000001111101111000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000001111101111000000000000};
            #100 x={28'b0000001111110001000000000000};
            #100 x={28'b0000001111110101000000000000};
            #100 x={28'b0000001111110101000000000000};
            #100 x={28'b0000001111110111000000000000};
            #100 x={28'b0000001111110110000000000000};
            #100 x={28'b0000001111110001000000000000};
            #100 x={28'b0000001111110101000000000000};
            #100 x={28'b0000001111111001000000000000};
            #100 x={28'b0000001111111001000000000000};
            #100 x={28'b0000001111111001000000000000};
            #100 x={28'b0000001111110110000000000000};
            #100 x={28'b0000001111110110000000000000};
            #100 x={28'b0000001111111000000000000000};
            #100 x={28'b0000001111111011000000000000};
            #100 x={28'b0000001111111010000000000000};
            #100 x={28'b0000001111111100000000000000};
            #100 x={28'b0000001111110111000000000000};
            #100 x={28'b0000001111110001000000000000};
            #100 x={28'b0000001111101101000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000001111110000000000000000};
            #100 x={28'b0000001111110000000000000000};
            #100 x={28'b0000001111101100000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111101100000000000000};
            #100 x={28'b0000001111110101000000000000};
            #100 x={28'b0000001111111010000000000000};
            #100 x={28'b0000001111110111000000000000};
            #100 x={28'b0000001111110001000000000000};
            #100 x={28'b0000001111110010000000000000};
            #100 x={28'b0000001111110100000000000000};
            #100 x={28'b0000001111110011000000000000};
            #100 x={28'b0000001111101111000000000000};
            #100 x={28'b0000001111101101000000000000};
            #100 x={28'b0000001111101101000000000000};
            #100 x={28'b0000001111101100000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000010000000011000000000000};
            #100 x={28'b0000010000101000000000000000};
            #100 x={28'b0000010001011001000000000000};
            #100 x={28'b0000010010010100000000000000};
            #100 x={28'b0000010011000011000000000000};
            #100 x={28'b0000010011001111000000000000};
            #100 x={28'b0000010010101110000000000000};
            #100 x={28'b0000010001110111000000000000};
            #100 x={28'b0000010001000100000000000000};
            #100 x={28'b0000010000011000000000000000};
            #100 x={28'b0000001111111000000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111101100000000000000};
            #100 x={28'b0000001111101100000000000000};
            #100 x={28'b0000001111101111000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000001111101101000000000000};
            #100 x={28'b0000001111101111000000000000};
            #100 x={28'b0000001111110010000000000000};
            #100 x={28'b0000001111111000000000000000};
            #100 x={28'b0000001111111000000000000000};
            #100 x={28'b0000001111110111000000000000};
            #100 x={28'b0000001111110110000000000000};
            #100 x={28'b0000001111110100000000000000};
            #100 x={28'b0000001111110100000000000000};
            #100 x={28'b0000001111111001000000000000};
            #100 x={28'b0000001111111100000000000000};
            #100 x={28'b0000001111111100000000000000};
            #100 x={28'b0000001111111000000000000000};
            #100 x={28'b0000001111110111000000000000};
            #100 x={28'b0000001111110101000000000000};
            #100 x={28'b0000001111110101000000000000};
            #100 x={28'b0000001111110101000000000000};
            #100 x={28'b0000001111110110000000000000};
            #100 x={28'b0000001111110100000000000000};
            #100 x={28'b0000001111110010000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111101101000000000000};
            #100 x={28'b0000001111110001000000000000};
            #100 x={28'b0000001111110001000000000000};
            #100 x={28'b0000001111101111000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000010000000101000000000000};
            #100 x={28'b0000010000110010000000000000};
            #100 x={28'b0000010001110000000000000000};
            #100 x={28'b0000010010110010000000000000};
            #100 x={28'b0000010011100101000000000000};
            #100 x={28'b0000010011100001000000000000};
            #100 x={28'b0000010010100111000000000000};
            #100 x={28'b0000010001100011000000000000};
            #100 x={28'b0000010000101000000000000000};
            #100 x={28'b0000010000000100000000000000};
            #100 x={28'b0000001111110101000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110011001000000000000};
            #100 x={28'b0000001110010100000000000000};
            #100 x={28'b0000001110010010000000000000};
            #100 x={28'b0000001110011010000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110010101000000000000};
            #100 x={28'b0000001110010010000000000000};
            #100 x={28'b0000001110001110000000000000};
            #100 x={28'b0000001110001110000000000000};
            #100 x={28'b0000001110010110000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000010000011111000000000000};
            #100 x={28'b0000010001100110000000000000};
            #100 x={28'b0000010010110000000000000000};
            #100 x={28'b0000010011100010000000000000};
            #100 x={28'b0000010011011100000000000000};
            #100 x={28'b0000010010101000000000000000};
            #100 x={28'b0000010001100011000000000000};
            #100 x={28'b0000010000011100000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110010010000000000000};
            #100 x={28'b0000001110001111000000000000};
            #100 x={28'b0000001110001101000000000000};
            #100 x={28'b0000001110000111000000000000};
            #100 x={28'b0000001110000110000000000000};
            #100 x={28'b0000001110000110000000000000};
            #100 x={28'b0000001110001101000000000000};
            #100 x={28'b0000001110010000000000000000};
            #100 x={28'b0000001110001100000000000000};
            #100 x={28'b0000001110001000000000000000};
            #100 x={28'b0000001110001000000000000000};
            #100 x={28'b0000001110000111000000000000};
            #100 x={28'b0000001110001100000000000000};
            #100 x={28'b0000001110001011000000000000};
            #100 x={28'b0000001110001001000000000000};
            #100 x={28'b0000001110000011000000000000};
            #100 x={28'b0000001110000001000000000000};
            #100 x={28'b0000001110000000000000000000};
            #100 x={28'b0000001110000010000000000000};
            #100 x={28'b0000001110001010000000000000};
            #100 x={28'b0000001110001111000000000000};
            #100 x={28'b0000001110001100000000000000};
            #100 x={28'b0000001110001000000000000000};
            #100 x={28'b0000001110000010000000000000};
            #100 x={28'b0000001110000001000000000000};
            #100 x={28'b0000001110000110000000000000};
            #100 x={28'b0000001110001001000000000000};
            #100 x={28'b0000001110000111000000000000};
            #100 x={28'b0000001110001001000000000000};
            #100 x={28'b0000001110001101000000000000};
            #100 x={28'b0000001110001100000000000000};
            #100 x={28'b0000001110000011000000000000};
            #100 x={28'b0000001101111100000000000000};
            #100 x={28'b0000001110000011000000000000};
            #100 x={28'b0000001110001011000000000000};
            #100 x={28'b0000001110001011000000000000};
            #100 x={28'b0000001110001011000000000000};
            #100 x={28'b0000001110001000000000000000};
            #100 x={28'b0000001110001000000000000000};
            #100 x={28'b0000001110000110000000000000};
            #100 x={28'b0000001110001101000000000000};
            #100 x={28'b0000001110001111000000000000};
            #100 x={28'b0000001110001100000000000000};
            #100 x={28'b0000001110001010000000000000};
            #100 x={28'b0000001110000111000000000000};
            #100 x={28'b0000001110001000000000000000};
            #100 x={28'b0000001110001001000000000000};
            #100 x={28'b0000001110001011000000000000};
            #100 x={28'b0000001110001010000000000000};
            #100 x={28'b0000001110000101000000000000};
            #100 x={28'b0000001110000110000000000000};
            #100 x={28'b0000001110001010000000000000};
            #100 x={28'b0000001110001101000000000000};
            #100 x={28'b0000001110001110000000000000};
            #100 x={28'b0000001110010000000000000000};
            #100 x={28'b0000001110010010000000000000};
            #100 x={28'b0000001110010110000000000000};
            #100 x={28'b0000001110010011000000000000};
            #100 x={28'b0000001110001111000000000000};
            #100 x={28'b0000001110001101000000000000};
            #100 x={28'b0000001110001111000000000000};
            #100 x={28'b0000001110010011000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110011001000000000000};
            #100 x={28'b0000001110011000000000000000};
            #100 x={28'b0000001110011010000000000000};
            #100 x={28'b0000001110011101000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110011001000000000000};
            #100 x={28'b0000001110010110000000000000};
            #100 x={28'b0000001110010111000000000000};
            #100 x={28'b0000001110010111000000000000};
            #100 x={28'b0000001110010101000000000000};
            #100 x={28'b0000001110011101000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110010010000000000000};
            #100 x={28'b0000001110001010000000000000};
            #100 x={28'b0000001110001101000000000000};
            #100 x={28'b0000001110010011000000000000};
            #100 x={28'b0000001110010110000000000000};
            #100 x={28'b0000001110011001000000000000};
            #100 x={28'b0000001110010011000000000000};
            #100 x={28'b0000001110001111000000000000};
            #100 x={28'b0000001110011000000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110011000000000000000};
            #100 x={28'b0000001110010001000000000000};
            #100 x={28'b0000001110001011000000000000};
            #100 x={28'b0000001110001110000000000000};
            #100 x={28'b0000001110010010000000000000};
            #100 x={28'b0000001110010101000000000000};
            #100 x={28'b0000001110010001000000000000};
            #100 x={28'b0000001110001011000000000000};
            #100 x={28'b0000001110000101000000000000};
            #100 x={28'b0000001110001001000000000000};
            #100 x={28'b0000001110010100000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110001010000000000000};
            #100 x={28'b0000001110000101000000000000};
            #100 x={28'b0000001110001101000000000000};
            #100 x={28'b0000001110010111000000000000};
            #100 x={28'b0000001110011001000000000000};
            #100 x={28'b0000001110010110000000000000};
            #100 x={28'b0000001110010010000000000000};
            #100 x={28'b0000001110010011000000000000};
            #100 x={28'b0000001110011001000000000000};
            #100 x={28'b0000001110010111000000000000};
            #100 x={28'b0000001110010110000000000000};
            #100 x={28'b0000001110010101000000000000};
            #100 x={28'b0000001110010011000000000000};
            #100 x={28'b0000001110010110000000000000};
            #100 x={28'b0000001110011010000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110011000000000000000};
            #100 x={28'b0000001110010101000000000000};
            #100 x={28'b0000001110010111000000000000};
            #100 x={28'b0000001110011000000000000000};
            #100 x={28'b0000001110010101000000000000};
            #100 x={28'b0000001110010111000000000000};
            #100 x={28'b0000001110011001000000000000};
            #100 x={28'b0000001110010110000000000000};
            #100 x={28'b0000001110010011000000000000};
            #100 x={28'b0000001110010010000000000000};
            #100 x={28'b0000001110001110000000000000};
            #100 x={28'b0000001110010011000000000000};
            #100 x={28'b0000001110011001000000000000};
            #100 x={28'b0000001110011001000000000000};
            #100 x={28'b0000001110011000000000000000};
            #100 x={28'b0000001110010100000000000000};
            #100 x={28'b0000001110001111000000000000};
            #100 x={28'b0000001110011000000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110010011000000000000};
            #100 x={28'b0000001110001010000000000000};
            #100 x={28'b0000001110001100000000000000};
            #100 x={28'b0000001110010101000000000000};
            #100 x={28'b0000001110011010000000000000};
            #100 x={28'b0000001110011000000000000000};
            #100 x={28'b0000001110010110000000000000};
            #100 x={28'b0000001110010101000000000000};
            #100 x={28'b0000001110010111000000000000};
            #100 x={28'b0000001110010110000000000000};
            #100 x={28'b0000001110010101000000000000};
            #100 x={28'b0000001110010010000000000000};
            #100 x={28'b0000001110010000000000000000};
            #100 x={28'b0000001110001111000000000000};
            #100 x={28'b0000001110010101000000000000};
            #100 x={28'b0000001110010101000000000000};
            #100 x={28'b0000001110010101000000000000};
            #100 x={28'b0000001110010110000000000000};
            #100 x={28'b0000001110011010000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011000000000000000};
            #100 x={28'b0000001110010100000000000000};
            #100 x={28'b0000001110010101000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110011001000000000000};
            #100 x={28'b0000001110010110000000000000};
            #100 x={28'b0000001110010100000000000000};
            #100 x={28'b0000001110010010000000000000};
            #100 x={28'b0000001110010101000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110010101000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011101000000000000};
            #100 x={28'b0000001110011001000000000000};
            #100 x={28'b0000001110011010000000000000};
            #100 x={28'b0000001110011000000000000000};
            #100 x={28'b0000001110010101000000000000};
            #100 x={28'b0000001110010001000000000000};
            #100 x={28'b0000001110010011000000000000};
            #100 x={28'b0000001110011000000000000000};
            #100 x={28'b0000001110011010000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110010101000000000000};
            #100 x={28'b0000001110010010000000000000};
            #100 x={28'b0000001110010010000000000000};
            #100 x={28'b0000001110010001000000000000};
            #100 x={28'b0000001110001110000000000000};
            #100 x={28'b0000001110000111000000000000};
            #100 x={28'b0000001110000010000000000000};
            #100 x={28'b0000001110000111000000000000};
            #100 x={28'b0000001110011101000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111111000000000000000};
            #100 x={28'b0000010000111001000000000000};
            #100 x={28'b0000010010000010000000000000};
            #100 x={28'b0000010011001100000000000000};
            #100 x={28'b0000010011111010000000000000};
            #100 x={28'b0000010011111001000000000000};
            #100 x={28'b0000010011000001000000000000};
            #100 x={28'b0000010001101010000000000000};
            #100 x={28'b0000010000100101000000000000};
            #100 x={28'b0000001111110111000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110010111000000000000};
            #100 x={28'b0000001110010100000000000000};
            #100 x={28'b0000001110011001000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110011010000000000000};
            #100 x={28'b0000001110010100000000000000};
            #100 x={28'b0000001110001110000000000000};
            #100 x={28'b0000001110001010000000000000};
            #100 x={28'b0000001110001001000000000000};
            #100 x={28'b0000001110010000000000000000};
            #100 x={28'b0000001110010001000000000000};
            #100 x={28'b0000001110010000000000000000};
            #100 x={28'b0000001110001110000000000000};
            #100 x={28'b0000001110010000000000000000};
            #100 x={28'b0000001110010010000000000000};
            #100 x={28'b0000001110010011000000000000};
            #100 x={28'b0000001110001111000000000000};
            #100 x={28'b0000001110001001000000000000};
            #100 x={28'b0000001110000110000000000000};
            #100 x={28'b0000001110001000000000000000};
            #100 x={28'b0000001110001110000000000000};
            #100 x={28'b0000001110010011000000000000};
            #100 x={28'b0000001110010011000000000000};
            #100 x={28'b0000001110010011000000000000};
            #100 x={28'b0000001110010100000000000000};
            #100 x={28'b0000001110011000000000000000};
            #100 x={28'b0000001110011010000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110011000000000000000};
            #100 x={28'b0000001110010100000000000000};
            #100 x={28'b0000001110010010000000000000};
            #100 x={28'b0000001110010001000000000000};
            #100 x={28'b0000001110010101000000000000};
            #100 x={28'b0000001110011000000000000000};
            #100 x={28'b0000001110011000000000000000};
            #100 x={28'b0000001110010101000000000000};
            #100 x={28'b0000001110010101000000000000};
            #100 x={28'b0000001110011001000000000000};
            #100 x={28'b0000001110010101000000000000};
            #100 x={28'b0000001110010010000000000000};
            #100 x={28'b0000001110001101000000000000};
            #100 x={28'b0000001110000101000000000000};
            #100 x={28'b0000001110001110000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110010111000000000000};
            #100 x={28'b0000001110011010000000000000};
            #100 x={28'b0000001110011010000000000000};
            #100 x={28'b0000001110011000000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110011001000000000000};
            #100 x={28'b0000001110010011000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111101100000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111110011000000000000};
            #100 x={28'b0000001111101011000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110010011000000000000};
            #100 x={28'b0000001110010010000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110011101000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110010101000000000000};
            #100 x={28'b0000001110011101000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110011001000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111101101000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110010101000000000000};
            #100 x={28'b0000001110001111000000000000};
            #100 x={28'b0000001110010001000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111110011000000000000};
            #100 x={28'b0000010000110010000000000000};
            #100 x={28'b0000010001111101000000000000};
            #100 x={28'b0000010011010001000000000000};
            #100 x={28'b0000010100010011000000000000};
            #100 x={28'b0000010100100011000000000000};
            #100 x={28'b0000010011110110000000000000};
            #100 x={28'b0000010010100101000000000000};
            #100 x={28'b0000010001010110000000000000};
            #100 x={28'b0000010000010111000000000000};
            #100 x={28'b0000010000000010000000000000};
            #100 x={28'b0000010000000011000000000000};
            #100 x={28'b0000001111101101000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110010101000000000000};
            #100 x={28'b0000001110011001000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110011101000000000000};
            #100 x={28'b0000001110010111000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110010110000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110011101000000000000};
            #100 x={28'b0000001110001101000000000000};
            #100 x={28'b0000001110001000000000000000};
            #100 x={28'b0000001110010001000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110011010000000000000};
            #100 x={28'b0000001110011010000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110011000000000000000};
            #100 x={28'b0000001110010010000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111101011000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111110001000000000000};
            #100 x={28'b0000001111111011000000000000};
            #100 x={28'b0000001111111000000000000000};
            #100 x={28'b0000001111110111000000000000};
            #100 x={28'b0000001111111001000000000000};
            #100 x={28'b0000001111110001000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111110110000000000000};
            #100 x={28'b0000001111111001000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111110001000000000000};
            #100 x={28'b0000010000100110000000000000};
            #100 x={28'b0000010001100011000000000000};
            #100 x={28'b0000010010101010000000000000};
            #100 x={28'b0000010011101111000000000000};
            #100 x={28'b0000010100011110000000000000};
            #100 x={28'b0000010100011100000000000000};
            #100 x={28'b0000010011101011000000000000};
            #100 x={28'b0000010010100100000000000000};
            #100 x={28'b0000010001011111000000000000};
            #100 x={28'b0000010000101111000000000000};
            #100 x={28'b0000010000011010000000000000};
            #100 x={28'b0000010000001000000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111101011000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000001111101101000000000000};
            #100 x={28'b0000001111110100000000000000};
            #100 x={28'b0000010000000000000000000000};
            #100 x={28'b0000001111111111000000000000};
            #100 x={28'b0000001111110011000000000000};
            #100 x={28'b0000001111101101000000000000};
            #100 x={28'b0000001111110000000000000000};
            #100 x={28'b0000001111111100000000000000};
            #100 x={28'b0000010000001000000000000000};
            #100 x={28'b0000010000001011000000000000};
            #100 x={28'b0000010000000100000000000000};
            #100 x={28'b0000001111111111000000000000};
            #100 x={28'b0000010000000000000000000000};
            #100 x={28'b0000001111111111000000000000};
            #100 x={28'b0000001111111110000000000000};
            #100 x={28'b0000001111111010000000000000};
            #100 x={28'b0000001111110011000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111101100000000000000};
            #100 x={28'b0000001111110011000000000000};
            #100 x={28'b0000001111101011000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111110110000000000000};
            #100 x={28'b0000001111111010000000000000};
            #100 x={28'b0000001111111101000000000000};
            #100 x={28'b0000001111110111000000000000};
            #100 x={28'b0000001111101111000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111110000000000000000};
            #100 x={28'b0000001111110011000000000000};
            #100 x={28'b0000001111110001000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111110011000000000000};
            #100 x={28'b0000001111110010000000000000};
            #100 x={28'b0000001111101100000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111110110000000000000};
            #100 x={28'b0000001111110000000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111110010000000000000};
            #100 x={28'b0000010000010111000000000000};
            #100 x={28'b0000010001001110000000000000};
            #100 x={28'b0000010010010011000000000000};
            #100 x={28'b0000010011011111000000000000};
            #100 x={28'b0000010100100000000000000000};
            #100 x={28'b0000010100111110000000000000};
            #100 x={28'b0000010100101101000000000000};
            #100 x={28'b0000010011101111000000000000};
            #100 x={28'b0000010010100101000000000000};
            #100 x={28'b0000010001100001000000000000};
            #100 x={28'b0000010000101011000000000000};
            #100 x={28'b0000010000011011000000000000};
            #100 x={28'b0000010000011010000000000000};
            #100 x={28'b0000010000001010000000000000};
            #100 x={28'b0000001111101011000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000001111110110000000000000};
            #100 x={28'b0000010000000000000000000000};
            #100 x={28'b0000010000000011000000000000};
            #100 x={28'b0000001111111100000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111110001000000000000};
            #100 x={28'b0000001111111110000000000000};
            #100 x={28'b0000010000000000000000000000};
            #100 x={28'b0000010000000001000000000000};
            #100 x={28'b0000010000000001000000000000};
            #100 x={28'b0000010000000001000000000000};
            #100 x={28'b0000010000000101000000000000};
            #100 x={28'b0000010000001111000000000000};
            #100 x={28'b0000010000001101000000000000};
            #100 x={28'b0000010000000011000000000000};
            #100 x={28'b0000001111111011000000000000};
            #100 x={28'b0000001111111100000000000000};
            #100 x={28'b0000010000000101000000000000};
            #100 x={28'b0000010000000111000000000000};
            #100 x={28'b0000010000000010000000000000};
            #100 x={28'b0000001111111001000000000000};
            #100 x={28'b0000001111110111000000000000};
            #100 x={28'b0000001111110100000000000000};
            #100 x={28'b0000001111110000000000000000};
            #100 x={28'b0000001111110001000000000000};
            #100 x={28'b0000001111101011000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111111011000000000000};
            #100 x={28'b0000010000000011000000000000};
            #100 x={28'b0000001111111100000000000000};
            #100 x={28'b0000001111110111000000000000};
            #100 x={28'b0000001111110010000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111110100000000000000};
            #100 x={28'b0000010000101110000000000000};
            #100 x={28'b0000010001101111000000000000};
            #100 x={28'b0000010010110110000000000000};
            #100 x={28'b0000010011111001000000000000};
            #100 x={28'b0000010100101001000000000000};
            #100 x={28'b0000010100101110000000000000};
            #100 x={28'b0000010100000000000000000000};
            #100 x={28'b0000010010110010000000000000};
            #100 x={28'b0000010001100100000000000000};
            #100 x={28'b0000010000100101000000000000};
            #100 x={28'b0000001111111010000000000000};
            #100 x={28'b0000001111101111000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000001111110011000000000000};
            #100 x={28'b0000001111110001000000000000};
            #100 x={28'b0000001111101100000000000000};
            #100 x={28'b0000001111101011000000000000};
            #100 x={28'b0000001111110010000000000000};
            #100 x={28'b0000001111110110000000000000};
            #100 x={28'b0000001111111000000000000000};
            #100 x={28'b0000001111111101000000000000};
            #100 x={28'b0000001111111010000000000000};
            #100 x={28'b0000001111110111000000000000};
            #100 x={28'b0000001111110100000000000000};
            #100 x={28'b0000001111111000000000000000};
            #100 x={28'b0000010000000001000000000000};
            #100 x={28'b0000010000000100000000000000};
            #100 x={28'b0000010000000010000000000000};
            #100 x={28'b0000001111111110000000000000};
            #100 x={28'b0000001111111100000000000000};
            #100 x={28'b0000001111111101000000000000};
            #100 x={28'b0000010000000011000000000000};
            #100 x={28'b0000010000000001000000000000};
            #100 x={28'b0000001111111101000000000000};
            #100 x={28'b0000001111110101000000000000};
            #100 x={28'b0000001111110011000000000000};
            #100 x={28'b0000001111110010000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111101111000000000000};
            #100 x={28'b0000001111110110000000000000};
            #100 x={28'b0000001111110111000000000000};
            #100 x={28'b0000001111110101000000000000};
            #100 x={28'b0000001111110001000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000001111101111000000000000};
            #100 x={28'b0000001111101101000000000000};
            #100 x={28'b0000001111110010000000000000};
            #100 x={28'b0000001111110000000000000000};
            #100 x={28'b0000001111101101000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111110000000000000000};
            #100 x={28'b0000010000011100000000000000};
            #100 x={28'b0000010001010011000000000000};
            #100 x={28'b0000010010010010000000000000};
            #100 x={28'b0000010011010111000000000000};
            #100 x={28'b0000010100010010000000000000};
            #100 x={28'b0000010100101011000000000000};
            #100 x={28'b0000010100010000000000000000};
            #100 x={28'b0000010011001101000000000000};
            #100 x={28'b0000010010000101000000000000};
            #100 x={28'b0000010000111111000000000000};
            #100 x={28'b0000010000001000000000000000};
            #100 x={28'b0000001111110011000000000000};
            #100 x={28'b0000001111110110000000000000};
            #100 x={28'b0000001111110001000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000001111110001000000000000};
            #100 x={28'b0000001111110011000000000000};
            #100 x={28'b0000001111110001000000000000};
            #100 x={28'b0000001111110010000000000000};
            #100 x={28'b0000001111110011000000000000};
            #100 x={28'b0000001111110111000000000000};
            #100 x={28'b0000001111111001000000000000};
            #100 x={28'b0000001111111000000000000000};
            #100 x={28'b0000001111110111000000000000};
            #100 x={28'b0000001111110011000000000000};
            #100 x={28'b0000001111110001000000000000};
            #100 x={28'b0000001111110001000000000000};
            #100 x={28'b0000001111110001000000000000};
            #100 x={28'b0000001111110001000000000000};
            #100 x={28'b0000001111101011000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111101011000000000000};
            #100 x={28'b0000001111101101000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000010000001101000000000000};
            #100 x={28'b0000010001000101000000000000};
            #100 x={28'b0000010010000011000000000000};
            #100 x={28'b0000010011001000000000000000};
            #100 x={28'b0000010100000011000000000000};
            #100 x={28'b0000010100001111000000000000};
            #100 x={28'b0000010011100001000000000000};
            #100 x={28'b0000010010010110000000000000};
            #100 x={28'b0000010001001100000000000000};
            #100 x={28'b0000010000001011000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110011101000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011101000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011101000000000000};
            #100 x={28'b0000001110011010000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111101011000000000000};
            #100 x={28'b0000001111101100000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111110001000000000000};
            #100 x={28'b0000010000100000000000000000};
            #100 x={28'b0000010001100010000000000000};
            #100 x={28'b0000010010100001000000000000};
            #100 x={28'b0000010011011110000000000000};
            #100 x={28'b0000010011111110000000000000};
            #100 x={28'b0000010011101011000000000000};
            #100 x={28'b0000010010101010000000000000};
            #100 x={28'b0000010001100001000000000000};
            #100 x={28'b0000010000101001000000000000};
            #100 x={28'b0000010000000000000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110011101000000000000};
            #100 x={28'b0000001110011010000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110011101000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110011101000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110011010000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110010111000000000000};
            #100 x={28'b0000001110011001000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110011000000000000000};
            #100 x={28'b0000001110010110000000000000};
            #100 x={28'b0000001110011000000000000000};
            #100 x={28'b0000001110011010000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110011001000000000000};
            #100 x={28'b0000001110011000000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110011101000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110011101000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110011010000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110010111000000000000};
            #100 x={28'b0000001110010101000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000010000010001000000000000};
            #100 x={28'b0000010001010101000000000000};
            #100 x={28'b0000010010011111000000000000};
            #100 x={28'b0000010011011110000000000000};
            #100 x={28'b0000010011110111000000000000};
            #100 x={28'b0000010011001111000000000000};
            #100 x={28'b0000010010000001000000000000};
            #100 x={28'b0000010000110110000000000000};
            #100 x={28'b0000001111111011000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110010101000000000000};
            #100 x={28'b0000001110010110000000000000};
            #100 x={28'b0000001110010111000000000000};
            #100 x={28'b0000001110011000000000000000};
            #100 x={28'b0000001110010010000000000000};
            #100 x={28'b0000001110010001000000000000};
            #100 x={28'b0000001110001111000000000000};
            #100 x={28'b0000001110010000000000000000};
            #100 x={28'b0000001110010110000000000000};
            #100 x={28'b0000001110011001000000000000};
            #100 x={28'b0000001110011000000000000000};
            #100 x={28'b0000001110010110000000000000};
            #100 x={28'b0000001110010011000000000000};
            #100 x={28'b0000001110010101000000000000};
            #100 x={28'b0000001110010111000000000000};
            #100 x={28'b0000001110010101000000000000};
            #100 x={28'b0000001110010011000000000000};
            #100 x={28'b0000001110010010000000000000};
            #100 x={28'b0000001110010000000000000000};
            #100 x={28'b0000001110010100000000000000};
            #100 x={28'b0000001110010110000000000000};
            #100 x={28'b0000001110011000000000000000};
            #100 x={28'b0000001110010110000000000000};
            #100 x={28'b0000001110010011000000000000};
            #100 x={28'b0000001110010010000000000000};
            #100 x={28'b0000001110010110000000000000};
            #100 x={28'b0000001110011000000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110011101000000000000};
            #100 x={28'b0000001110011010000000000000};
            #100 x={28'b0000001110010101000000000000};
            #100 x={28'b0000001110010011000000000000};
            #100 x={28'b0000001110011001000000000000};
            #100 x={28'b0000001110011010000000000000};
            #100 x={28'b0000001110011001000000000000};
            #100 x={28'b0000001110011010000000000000};
            #100 x={28'b0000001110011010000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110011010000000000000};
            #100 x={28'b0000001110011010000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110011010000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111101011000000000000};
            #100 x={28'b0000001111101100000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000010000010110000000000000};
            #100 x={28'b0000010001001110000000000000};
            #100 x={28'b0000010010000111000000000000};
            #100 x={28'b0000010011010010000000000000};
            #100 x={28'b0000010100010001000000000000};
            #100 x={28'b0000010100011001000000000000};
            #100 x={28'b0000010011100010000000000000};
            #100 x={28'b0000010010011011000000000000};
            #100 x={28'b0000010001010111000000000000};
            #100 x={28'b0000010000010011000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110010000000000000000};
            #100 x={28'b0000001110010100000000000000};
            #100 x={28'b0000001110011101000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110010111000000000000};
            #100 x={28'b0000001110010011000000000000};
            #100 x={28'b0000001110011000000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110010101000000000000};
            #100 x={28'b0000001110001101000000000000};
            #100 x={28'b0000001110010110000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110011010000000000000};
            #100 x={28'b0000001110010100000000000000};
            #100 x={28'b0000001110010010000000000000};
            #100 x={28'b0000001110011001000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110011101000000000000};
            #100 x={28'b0000001110001100000000000000};
            #100 x={28'b0000001110000100000000000000};
            #100 x={28'b0000001110000110000000000000};
            #100 x={28'b0000001110001111000000000000};
            #100 x={28'b0000001110011101000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110011010000000000000};
            #100 x={28'b0000001110001000000000000000};
            #100 x={28'b0000001110000100000000000000};
            #100 x={28'b0000001110001111000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110011001000000000000};
            #100 x={28'b0000001110011000000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110011010000000000000};
            #100 x={28'b0000001110010101000000000000};
            #100 x={28'b0000001110011000000000000000};
            #100 x={28'b0000001110010101000000000000};
            #100 x={28'b0000001110010010000000000000};
            #100 x={28'b0000001110010000000000000000};
            #100 x={28'b0000001110010100000000000000};
            #100 x={28'b0000001110011010000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011011000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110010111000000000000};
            #100 x={28'b0000001110011000000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011101000000000000};
            #100 x={28'b0000001110011100000000000000};
            #100 x={28'b0000001110011101000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111101101000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000010000000100000000000000};
            #100 x={28'b0000010000110100000000000000};
            #100 x={28'b0000010001110110000000000000};
            #100 x={28'b0000010010111111000000000000};
            #100 x={28'b0000010100001001000000000000};
            #100 x={28'b0000010100101101000000000000};
            #100 x={28'b0000010100011001000000000000};
            #100 x={28'b0000010011010101000000000000};
            #100 x={28'b0000010010001101000000000000};
            #100 x={28'b0000010001001101000000000000};
            #100 x={28'b0000010000100010000000000000};
            #100 x={28'b0000010000001110000000000000};
            #100 x={28'b0000010000001011000000000000};
            #100 x={28'b0000001111111111000000000000};
            #100 x={28'b0000001111110010000000000000};
            #100 x={28'b0000001111110001000000000000};
            #100 x={28'b0000001111101101000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111101100000000000000};
            #100 x={28'b0000001111110010000000000000};
            #100 x={28'b0000001111110011000000000000};
            #100 x={28'b0000001111110001000000000000};
            #100 x={28'b0000001111110011000000000000};
            #100 x={28'b0000001111111001000000000000};
            #100 x={28'b0000010000000001000000000000};
            #100 x={28'b0000010000000001000000000000};
            #100 x={28'b0000001111111011000000000000};
            #100 x={28'b0000001111111010000000000000};
            #100 x={28'b0000010000000000000000000000};
            #100 x={28'b0000010000000011000000000000};
            #100 x={28'b0000010000001001000000000000};
            #100 x={28'b0000010000000110000000000000};
            #100 x={28'b0000010000000101000000000000};
            #100 x={28'b0000010000000101000000000000};
            #100 x={28'b0000010000000111000000000000};
            #100 x={28'b0000010000000110000000000000};
            #100 x={28'b0000010000000111000000000000};
            #100 x={28'b0000010000000101000000000000};
            #100 x={28'b0000010000000011000000000000};
            #100 x={28'b0000001111111111000000000000};
            #100 x={28'b0000001111111010000000000000};
            #100 x={28'b0000001111111011000000000000};
            #100 x={28'b0000001111111101000000000000};
            #100 x={28'b0000001111111011000000000000};
            #100 x={28'b0000001111110111000000000000};
            #100 x={28'b0000001111110101000000000000};
            #100 x={28'b0000001111110011000000000000};
            #100 x={28'b0000001111101111000000000000};
            #100 x={28'b0000001111101100000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111101011000000000000};
            #100 x={28'b0000001111110000000000000000};
            #100 x={28'b0000001111110110000000000000};
            #100 x={28'b0000001111110100000000000000};
            #100 x={28'b0000001111110000000000000000};
            #100 x={28'b0000001111110010000000000000};
            #100 x={28'b0000001111110111000000000000};
            #100 x={28'b0000001111111100000000000000};
            #100 x={28'b0000010000000010000000000000};
            #100 x={28'b0000010000000110000000000000};
            #100 x={28'b0000010000001101000000000000};
            #100 x={28'b0000010000010000000000000000};
            #100 x={28'b0000010000010000000000000000};
            #100 x={28'b0000010000001101000000000000};
            #100 x={28'b0000010000001010000000000000};
            #100 x={28'b0000010000001001000000000000};
            #100 x={28'b0000010000000111000000000000};
            #100 x={28'b0000010000000110000000000000};
            #100 x={28'b0000010000000110000000000000};
            #100 x={28'b0000010000000110000000000000};
            #100 x={28'b0000010000000110000000000000};
            #100 x={28'b0000010000000100000000000000};
            #100 x={28'b0000001111111110000000000000};
            #100 x={28'b0000001111111100000000000000};
            #100 x={28'b0000001111111011000000000000};
            #100 x={28'b0000001111111011000000000000};
            #100 x={28'b0000001111110111000000000000};
            #100 x={28'b0000001111110100000000000000};
            #100 x={28'b0000001111110010000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111110000000000000000};
            #100 x={28'b0000010000010111000000000000};
            #100 x={28'b0000010001000100000000000000};
            #100 x={28'b0000010001111000000000000000};
            #100 x={28'b0000010010111001000000000000};
            #100 x={28'b0000010011111110000000000000};
            #100 x={28'b0000010100101110000000000000};
            #100 x={28'b0000010100101111000000000000};
            #100 x={28'b0000010011111011000000000000};
            #100 x={28'b0000010010110110000000000000};
            #100 x={28'b0000010001110100000000000000};
            #100 x={28'b0000010000111010000000000000};
            #100 x={28'b0000010000010111000000000000};
            #100 x={28'b0000010000010001000000000000};
            #100 x={28'b0000010000010011000000000000};
            #100 x={28'b0000010000001010000000000000};
            #100 x={28'b0000001111111001000000000000};
            #100 x={28'b0000001111110010000000000000};
            #100 x={28'b0000001111101111000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111101011000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111101100000000000000};
            #100 x={28'b0000001111110001000000000000};
            #100 x={28'b0000001111110111000000000000};
            #100 x={28'b0000001111111000000000000000};
            #100 x={28'b0000001111111001000000000000};
            #100 x={28'b0000001111111000000000000000};
            #100 x={28'b0000001111111100000000000000};
            #100 x={28'b0000010000000000000000000000};
            #100 x={28'b0000010000000000000000000000};
            #100 x={28'b0000010000000000000000000000};
            #100 x={28'b0000010000000001000000000000};
            #100 x={28'b0000010000000011000000000000};
            #100 x={28'b0000010000000110000000000000};
            #100 x={28'b0000010000000111000000000000};
            #100 x={28'b0000010000001011000000000000};
            #100 x={28'b0000010000000111000000000000};
            #100 x={28'b0000010000001101000000000000};
            #100 x={28'b0000010000001100000000000000};
            #100 x={28'b0000010000001010000000000000};
            #100 x={28'b0000010000001001000000000000};
            #100 x={28'b0000010000001011000000000000};
            #100 x={28'b0000010000001101000000000000};
            #100 x={28'b0000010000001101000000000000};
            #100 x={28'b0000010000001001000000000000};
            #100 x={28'b0000010000000011000000000000};
            #100 x={28'b0000001111111111000000000000};
            #100 x={28'b0000001111111101000000000000};
            #100 x={28'b0000001111111100000000000000};
            #100 x={28'b0000001111111000000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000001111101011000000000000};
            #100 x={28'b0000001111101111000000000000};
            #100 x={28'b0000001111110001000000000000};
            #100 x={28'b0000001111101101000000000000};
            #100 x={28'b0000001111101100000000000000};
            #100 x={28'b0000001111101100000000000000};
            #100 x={28'b0000001111101011000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111101111000000000000};
            #100 x={28'b0000001111110011000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111110101000000000000};
            #100 x={28'b0000010000000000000000000000};
            #100 x={28'b0000010000000000000000000000};
            #100 x={28'b0000001111110111000000000000};
            #100 x={28'b0000001111101111000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111101100000000000000};
            #100 x={28'b0000001111110001000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000010000010010000000000000};
            #100 x={28'b0000010001000011000000000000};
            #100 x={28'b0000010001111110000000000000};
            #100 x={28'b0000010011000110000000000000};
            #100 x={28'b0000010100001001000000000000};
            #100 x={28'b0000010100100111000000000000};
            #100 x={28'b0000010100001011000000000000};
            #100 x={28'b0000010011001111000000000000};
            #100 x={28'b0000010010001111000000000000};
            #100 x={28'b0000010001010100000000000000};
            #100 x={28'b0000010000101001000000000000};
            #100 x={28'b0000010000001110000000000000};
            #100 x={28'b0000010000001010000000000000};
            #100 x={28'b0000010000000101000000000000};
            #100 x={28'b0000001111111101000000000000};
            #100 x={28'b0000001111111000000000000000};
            #100 x={28'b0000001111111010000000000000};
            #100 x={28'b0000001111111000000000000000};
            #100 x={28'b0000001111101101000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111110001000000000000};
            #100 x={28'b0000001111111000000000000000};
            #100 x={28'b0000001111110101000000000000};
            #100 x={28'b0000001111110011000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000010000000100000000000000};
            #100 x={28'b0000010000010111000000000000};
            #100 x={28'b0000010000010100000000000000};
            #100 x={28'b0000010000000101000000000000};
            #100 x={28'b0000001111101100000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111111000000000000000};
            #100 x={28'b0000001111111001000000000000};
            #100 x={28'b0000001111101011000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111110001000000000000};
            #100 x={28'b0000010000010111000000000000};
            #100 x={28'b0000010000101011000000000000};
            #100 x={28'b0000010000010101000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000010000011111000000000000};
            #100 x={28'b0000010000110010000000000000};
            #100 x={28'b0000010000011110000000000000};
            #100 x={28'b0000001111111000000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111101011000000000000};
            #100 x={28'b0000001111110010000000000000};
            #100 x={28'b0000010000000111000000000000};
            #100 x={28'b0000010000101011000000000000};
            #100 x={28'b0000010001000110000000000000};
            #100 x={28'b0000010000111110000000000000};
            #100 x={28'b0000010000011100000000000000};
            #100 x={28'b0000001111110101000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000010000010100000000000000};
            #100 x={28'b0000010001000100000000000000};
            #100 x={28'b0000010001011100000000000000};
            #100 x={28'b0000010001010100000000000000};
            #100 x={28'b0000010000110111000000000000};
            #100 x={28'b0000010000001110000000000000};
            #100 x={28'b0000001111110001000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000010000000100000000000000};
            #100 x={28'b0000010000011110000000000000};
            #100 x={28'b0000010000101000000000000000};
            #100 x={28'b0000010000100101000000000000};
            #100 x={28'b0000010000011010000000000000};
            #100 x={28'b0000010000000101000000000000};
            #100 x={28'b0000001111110110000000000000};
            #100 x={28'b0000001111111001000000000000};
            #100 x={28'b0000010000010000000000000000};
            #100 x={28'b0000010000101010000000000000};
            #100 x={28'b0000010000101011000000000000};
            #100 x={28'b0000010000010000000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111110110000000000000};
            #100 x={28'b0000001111111100000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111111101000000000000};
            #100 x={28'b0000010000001100000000000000};
            #100 x={28'b0000010000001001000000000000};
            #100 x={28'b0000010000000101000000000000};
            #100 x={28'b0000001111111011000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111111011000000000000};
            #100 x={28'b0000010000001000000000000000};
            #100 x={28'b0000001111111110000000000000};
            #100 x={28'b0000001111101100000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111110000000000000000};
            #100 x={28'b0000001111110111000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111110001000000000000};
            #100 x={28'b0000001111111111000000000000};
            #100 x={28'b0000001111101100000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111101011000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111101111000000000000};
            #100 x={28'b0000001111111011000000000000};
            #100 x={28'b0000001111111100000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111101111000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111101111000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000001111101111000000000000};
            #100 x={28'b0000001111101111000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000001111101011000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111110110000000000000};
            #100 x={28'b0000010000100010000000000000};
            #100 x={28'b0000010001011101000000000000};
            #100 x={28'b0000010010100100000000000000};
            #100 x={28'b0000010011100100000000000000};
            #100 x={28'b0000010100000110000000000000};
            #100 x={28'b0000010011110001000000000000};
            #100 x={28'b0000010010110100000000000000};
            #100 x={28'b0000010001101111000000000000};
            #100 x={28'b0000010000111111000000000000};
            #100 x={28'b0000010000011101000000000000};
            #100 x={28'b0000010000001000000000000000};
            #100 x={28'b0000001111110110000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111101111000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000001111101100000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111101100000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000001111101101000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111110010000000000000};
            #100 x={28'b0000010000101000000000000000};
            #100 x={28'b0000010001100011000000000000};
            #100 x={28'b0000010010101010000000000000};
            #100 x={28'b0000010011100010000000000000};
            #100 x={28'b0000010011110111000000000000};
            #100 x={28'b0000010011011010000000000000};
            #100 x={28'b0000010010011101000000000000};
            #100 x={28'b0000010001100000000000000000};
            #100 x={28'b0000010000101101000000000000};
            #100 x={28'b0000010000000100000000000000};
            #100 x={28'b0000001111101111000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111101100000000000000};
            #100 x={28'b0000001111101011000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111101111000000000000};
            #100 x={28'b0000010000100000000000000000};
            #100 x={28'b0000010001010011000000000000};
            #100 x={28'b0000010010001111000000000000};
            #100 x={28'b0000010011001000000000000000};
            #100 x={28'b0000010011110000000000000000};
            #100 x={28'b0000010011101100000000000000};
            #100 x={28'b0000010010111000000000000000};
            #100 x={28'b0000010001111110000000000000};
            #100 x={28'b0000010001001010000000000000};
            #100 x={28'b0000010000011101000000000000};
            #100 x={28'b0000001111111101000000000000};
            #100 x={28'b0000001111110000000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111101101000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111101011000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000001111110000000000000000};
            #100 x={28'b0000001111101111000000000000};
            #100 x={28'b0000001111101101000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111101100000000000000};
            #100 x={28'b0000001111101100000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111101011000000000000};
            #100 x={28'b0000001111101011000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111110110000000000000};
            #100 x={28'b0000010000100110000000000000};
            #100 x={28'b0000010001011011000000000000};
            #100 x={28'b0000010010011011000000000000};
            #100 x={28'b0000010011010101000000000000};
            #100 x={28'b0000010011110011000000000000};
            #100 x={28'b0000010011011101000000000000};
            #100 x={28'b0000010010100011000000000000};
            #100 x={28'b0000010001100111000000000000};
            #100 x={28'b0000010000110011000000000000};
            #100 x={28'b0000010000000111000000000000};
            #100 x={28'b0000001111110101000000000000};
            #100 x={28'b0000001111110000000000000000};
            #100 x={28'b0000001111101011000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111101011000000000000};
            #100 x={28'b0000001111101100000000000000};
            #100 x={28'b0000001111101101000000000000};
            #100 x={28'b0000001111101101000000000000};
            #100 x={28'b0000001111101100000000000000};
            #100 x={28'b0000001111101101000000000000};
            #100 x={28'b0000001111101011000000000000};
            #100 x={28'b0000001111101111000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000001111101011000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111101100000000000000};
            #100 x={28'b0000010000010110000000000000};
            #100 x={28'b0000010001001011000000000000};
            #100 x={28'b0000010010001101000000000000};
            #100 x={28'b0000010011000111000000000000};
            #100 x={28'b0000010011011111000000000000};
            #100 x={28'b0000010011000101000000000000};
            #100 x={28'b0000010010001010000000000000};
            #100 x={28'b0000010001001101000000000000};
            #100 x={28'b0000010000011111000000000000};
            #100 x={28'b0000001111111110000000000000};
            #100 x={28'b0000001111101101000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110101000000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100000000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110011110000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100101000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100010000000000000};
            #100 x={28'b0000001110011111000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100100000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100001000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100011000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110100111000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110100110000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111110000000000000000};
            #100 x={28'b0000010000011010000000000000};
            #100 x={28'b0000010001000111000000000000};
            #100 x={28'b0000010001111100000000000000};
            #100 x={28'b0000010010110100000000000000};
            #100 x={28'b0000010011011101000000000000};
            #100 x={28'b0000010011011011000000000000};
            #100 x={28'b0000010010110001000000000000};
            #100 x={28'b0000010001111101000000000000};
            #100 x={28'b0000010001001101000000000000};
            #100 x={28'b0000010000100101000000000000};
            #100 x={28'b0000010000000100000000000000};
            #100 x={28'b0000001111110110000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111101011000000000000};
            #100 x={28'b0000001111101101000000000000};
            #100 x={28'b0000001111101101000000000000};
            #100 x={28'b0000001111101100000000000000};
            #100 x={28'b0000001111101101000000000000};
            #100 x={28'b0000001111110010000000000000};
            #100 x={28'b0000001111110100000000000000};
            #100 x={28'b0000001111110011000000000000};
            #100 x={28'b0000001111110001000000000000};
            #100 x={28'b0000001111110001000000000000};
            #100 x={28'b0000001111101100000000000000};
            #100 x={28'b0000001111101100000000000000};
            #100 x={28'b0000001111101101000000000000};
            #100 x={28'b0000001111101100000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111101100000000000000};
            #100 x={28'b0000001111110011000000000000};
            #100 x={28'b0000001111110111000000000000};
            #100 x={28'b0000001111111110000000000000};
            #100 x={28'b0000010000000000000000000000};
            #100 x={28'b0000010000000011000000000000};
            #100 x={28'b0000010000000011000000000000};
            #100 x={28'b0000010000000000000000000000};
            #100 x={28'b0000001111111110000000000000};
            #100 x={28'b0000001111111101000000000000};
            #100 x={28'b0000001111111001000000000000};
            #100 x={28'b0000001111110110000000000000};
            #100 x={28'b0000001111110111000000000000};
            #100 x={28'b0000001111110111000000000000};
            #100 x={28'b0000001111110110000000000000};
            #100 x={28'b0000001111110011000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000001111110000000000000000};
            #100 x={28'b0000001111110010000000000000};
            #100 x={28'b0000001111110010000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000010000001010000000000000};
            #100 x={28'b0000010000110011000000000000};
            #100 x={28'b0000010001100011000000000000};
            #100 x={28'b0000010010011000000000000000};
            #100 x={28'b0000010011001111000000000000};
            #100 x={28'b0000010011110101000000000000};
            #100 x={28'b0000010011111011000000000000};
            #100 x={28'b0000010011011001000000000000};
            #100 x={28'b0000010010100111000000000000};
            #100 x={28'b0000010001110110000000000000};
            #100 x={28'b0000010001001010000000000000};
            #100 x={28'b0000010000100101000000000000};
            #100 x={28'b0000010000010101000000000000};
            #100 x={28'b0000010000001100000000000000};
            #100 x={28'b0000010000000001000000000000};
            #100 x={28'b0000001111110100000000000000};
            #100 x={28'b0000001111110101000000000000};
            #100 x={28'b0000001111110010000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000001111101011000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111101100000000000000};
            #100 x={28'b0000001111110010000000000000};
            #100 x={28'b0000001111110101000000000000};
            #100 x={28'b0000001111111000000000000000};
            #100 x={28'b0000001111110110000000000000};
            #100 x={28'b0000001111110110000000000000};
            #100 x={28'b0000001111111000000000000000};
            #100 x={28'b0000001111111100000000000000};
            #100 x={28'b0000010000000000000000000000};
            #100 x={28'b0000010000000000000000000000};
            #100 x={28'b0000010000000001000000000000};
            #100 x={28'b0000010000000000000000000000};
            #100 x={28'b0000010000000100000000000000};
            #100 x={28'b0000010000000110000000000000};
            #100 x={28'b0000010000000111000000000000};
            #100 x={28'b0000010000000010000000000000};
            #100 x={28'b0000010000000101000000000000};
            #100 x={28'b0000010000000110000000000000};
            #100 x={28'b0000010000001001000000000000};
            #100 x={28'b0000010000001100000000000000};
            #100 x={28'b0000010000001100000000000000};
            #100 x={28'b0000010000001100000000000000};
            #100 x={28'b0000010000000111000000000000};
            #100 x={28'b0000010000001000000000000000};
            #100 x={28'b0000010000001001000000000000};
            #100 x={28'b0000010000001001000000000000};
            #100 x={28'b0000010000000111000000000000};
            #100 x={28'b0000010000000011000000000000};
            #100 x={28'b0000001111111111000000000000};
            #100 x={28'b0000001111111011000000000000};
            #100 x={28'b0000001111111010000000000000};
            #100 x={28'b0000001111111100000000000000};
            #100 x={28'b0000001111110110000000000000};
            #100 x={28'b0000001111110011000000000000};
            #100 x={28'b0000001111110011000000000000};
            #100 x={28'b0000001111110000000000000000};
            #100 x={28'b0000001111110001000000000000};
            #100 x={28'b0000001111101111000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111101011000000000000};
            #100 x={28'b0000001111101100000000000000};
            #100 x={28'b0000001111101100000000000000};
            #100 x={28'b0000001111101101000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111101110000000000000};
            #100 x={28'b0000001111110010000000000000};
            #100 x={28'b0000001111110111000000000000};
            #100 x={28'b0000001111111010000000000000};
            #100 x={28'b0000001111111011000000000000};
            #100 x={28'b0000010000000010000000000000};
            #100 x={28'b0000010000000011000000000000};
            #100 x={28'b0000010000001000000000000000};
            #100 x={28'b0000010000000110000000000000};
            #100 x={28'b0000010000000010000000000000};
            #100 x={28'b0000001111111111000000000000};
            #100 x={28'b0000001111111110000000000000};
            #100 x={28'b0000010000000000000000000000};
            #100 x={28'b0000001111111111000000000000};
            #100 x={28'b0000001111111101000000000000};
            #100 x={28'b0000001111111100000000000000};
            #100 x={28'b0000001111111000000000000000};
            #100 x={28'b0000001111110100000000000000};
            #100 x={28'b0000001111110100000000000000};
            #100 x={28'b0000001111110011000000000000};
            #100 x={28'b0000001111110010000000000000};
            #100 x={28'b0000001111101101000000000000};
            #100 x={28'b0000001111101011000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111110100000000000000};
            #100 x={28'b0000010000011000000000000000};
            #100 x={28'b0000010001000001000000000000};
            #100 x={28'b0000010001110011000000000000};
            #100 x={28'b0000010010101111000000000000};
            #100 x={28'b0000010011100100000000000000};
            #100 x={28'b0000010011110101000000000000};
            #100 x={28'b0000010011011110000000000000};
            #100 x={28'b0000010010100111000000000000};
            #100 x={28'b0000010001110100000000000000};
            #100 x={28'b0000010001000110000000000000};
            #100 x={28'b0000010000100100000000000000};
            #100 x={28'b0000010000010000000000000000};
            #100 x={28'b0000010000001101000000000000};
            #100 x={28'b0000010000000101000000000000};
            #100 x={28'b0000001111111011000000000000};
            #100 x={28'b0000001111110010000000000000};
            #100 x={28'b0000001111110010000000000000};
            #100 x={28'b0000001111101101000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111101101000000000000};
            #100 x={28'b0000001111110001000000000000};
            #100 x={28'b0000001111110010000000000000};
            #100 x={28'b0000001111110010000000000000};
            #100 x={28'b0000001111110011000000000000};
            #100 x={28'b0000001111110011000000000000};
            #100 x={28'b0000001111110111000000000000};
            #100 x={28'b0000001111111001000000000000};
            #100 x={28'b0000001111111011000000000000};
            #100 x={28'b0000001111111101000000000000};
            #100 x={28'b0000001111111101000000000000};
            #100 x={28'b0000001111111101000000000000};
            #100 x={28'b0000001111111100000000000000};
            #100 x={28'b0000001111111110000000000000};
            #100 x={28'b0000001111111111000000000000};
            #100 x={28'b0000010000000010000000000000};
            #100 x={28'b0000010000000000000000000000};
            #100 x={28'b0000001111111110000000000000};
            #100 x={28'b0000001111111110000000000000};
            #100 x={28'b0000001111111101000000000000};
            #100 x={28'b0000001111111011000000000000};
            #100 x={28'b0000001111111100000000000000};
            #100 x={28'b0000001111111010000000000000};
            #100 x={28'b0000001111110110000000000000};
            #100 x={28'b0000001111110011000000000000};
            #100 x={28'b0000001111110001000000000000};
            #100 x={28'b0000001111110001000000000000};
            #100 x={28'b0000001111101111000000000000};
            #100 x={28'b0000001111101011000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111110011000000000000};
            #100 x={28'b0000001111111000000000000000};
            #100 x={28'b0000001111111000000000000000};
            #100 x={28'b0000001111110110000000000000};
            #100 x={28'b0000001111110010000000000000};
            #100 x={28'b0000001111110010000000000000};
            #100 x={28'b0000001111110001000000000000};
            #100 x={28'b0000001111110110000000000000};
            #100 x={28'b0000001111110001000000000000};
            #100 x={28'b0000001111101101000000000000};
            #100 x={28'b0000001111101011000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000010000000001000000000000};
            #100 x={28'b0000010000101011000000000000};
            #100 x={28'b0000010001011011000000000000};
            #100 x={28'b0000010010010111000000000000};
            #100 x={28'b0000010011001010000000000000};
            #100 x={28'b0000010011010111000000000000};
            #100 x={28'b0000010010110110000000000000};
            #100 x={28'b0000010001111101000000000000};
            #100 x={28'b0000010001001000000000000000};
            #100 x={28'b0000010000100000000000000000};
            #100 x={28'b0000010000000111000000000000};
            #100 x={28'b0000001111111111000000000000};
            #100 x={28'b0000001111110111000000000000};
            #100 x={28'b0000001111101011000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111101011000000000000};
            #100 x={28'b0000001111101111000000000000};
            #100 x={28'b0000001111101100000000000000};
            #100 x={28'b0000001111101100000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111101011000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111111001000000000000};
            #100 x={28'b0000010000101011000000000000};
            #100 x={28'b0000010001100001000000000000};
            #100 x={28'b0000010010011101000000000000};
            #100 x={28'b0000010011001101000000000000};
            #100 x={28'b0000010011001011000000000000};
            #100 x={28'b0000010010011111000000000000};
            #100 x={28'b0000010001100101000000000000};
            #100 x={28'b0000010000110000000000000000};
            #100 x={28'b0000010000001010000000000000};
            #100 x={28'b0000001111111000000000000000};
            #100 x={28'b0000001111101101000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110011000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110110111000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111010010000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111101011000000000000};
            #100 x={28'b0000001111100111000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111101101000000000000};
            #100 x={28'b0000001111110000000000000000};
            #100 x={28'b0000001111110000000000000000};
            #100 x={28'b0000001111101101000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011100000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000101000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001010000000000000};
            #100 x={28'b0000001111001100000000000000};
            #100 x={28'b0000001111001110000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001011000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111011101000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111101010000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100001000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011011000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011000000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110110100000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000010000000011000000000000};
            #100 x={28'b0000010000110111000000000000};
            #100 x={28'b0000010001110000000000000000};
            #100 x={28'b0000010010101001000000000000};
            #100 x={28'b0000010011001101000000000000};
            #100 x={28'b0000010011000101000000000000};
            #100 x={28'b0000010010010100000000000000};
            #100 x={28'b0000010001011100000000000000};
            #100 x={28'b0000010000100110000000000000};
            #100 x={28'b0000010000000000000000000000};
            #100 x={28'b0000001111101111000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111000111000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101010000000000000};
            #100 x={28'b0000001110101001000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101100000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110101110000000000000};
            #100 x={28'b0000001110101101000000000000};
            #100 x={28'b0000001110101011000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110101000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110101111000000000000};
            #100 x={28'b0000001110110010000000000000};
            #100 x={28'b0000001110110001000000000000};
            #100 x={28'b0000001110110000000000000000};
            #100 x={28'b0000001110110110000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001000000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111001101000000000000};
            #100 x={28'b0000001111010000000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010101000000000000};
            #100 x={28'b0000001111010111000000000000};
            #100 x={28'b0000001111011010000000000000};
            #100 x={28'b0000001111011110000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111100101000000000000};
            #100 x={28'b0000001111100010000000000000};
            #100 x={28'b0000001111100100000000000000};
            #100 x={28'b0000001111101000000000000000};
            #100 x={28'b0000001111101100000000000000};
            #100 x={28'b0000001111101001000000000000};
            #100 x={28'b0000001111100110000000000000};
            #100 x={28'b0000001111100011000000000000};
            #100 x={28'b0000001111100000000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011111000000000000};
            #100 x={28'b0000001111011001000000000000};
            #100 x={28'b0000001111010110000000000000};
            #100 x={28'b0000001111010100000000000000};
            #100 x={28'b0000001111010011000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111010001000000000000};
            #100 x={28'b0000001111001111000000000000};
            #100 x={28'b0000001111001001000000000000};
            #100 x={28'b0000001111000110000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000100000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111011000000000000};
            #100 x={28'b0000001110111001000000000000};
            #100 x={28'b0000001110111010000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001110111100000000000000};
            #100 x={28'b0000001110111000000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111111000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000011000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001110111110000000000000};
            #100 x={28'b0000001110111101000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000010000000000000};
            #100 x={28'b0000001111000001000000000000};
            #100 x={28'b0000001111000000000000000000};
            #100 x={28'b0000001110111111000000000000};




        $finish;
    end

    // initial begin
    //      $monitor($time," x=%d y=%d",x,y);
    // end

    // initial begin
    //      $monitor(" x=%d",x);
    // end

    initial begin
         $monitor(" y=%d",y);
    end

    // Generate wave file
    initial begin
	$fsdbDumpfile("tb_pli.fsdb");
	$fsdbDumpvars;
	//$fsdbDumpMDA;
    end
      
endmodule